work.shiftr(main) rtlc_no_parameters
