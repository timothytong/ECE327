// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II"
// VERSION "Version 9.0 Build 132 02/25/2009 SJ Full Version"

// DATE "01/26/2016 18:37:17"

// 
// Device: Altera EP2C35F672C7 Package FBGA672
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module fir_top_chip (	clock_50,
	clock_27,
	key,
	sw,
	ledg,
	ledr,
	hex0,
	hex1,
	hex2,
	hex3,
	hex4,
	hex5,
	hex6,
	hex7,
	aud_xck,
	aud_bclk,
	aud_dacdat,
	aud_daclrck,
	aud_adclrck,
	i2c_sdat,
	i2c_sclk);
input 	clock_50;
input 	clock_27;
input 	[3:0] key;
input 	[17:0] sw;
output 	[8:0] ledg;
output 	[17:0] ledr;
output 	[6:0] hex0;
output 	[6:0] hex1;
output 	[6:0] hex2;
output 	[6:0] hex3;
output 	[6:0] hex4;
output 	[6:0] hex5;
output 	[6:0] hex6;
output 	[6:0] hex7;
output 	aud_xck;
inout 	aud_bclk;
output 	aud_dacdat;
output 	aud_daclrck;
output 	aud_adclrck;
inout 	i2c_sdat;
output 	i2c_sclk;

wire gnd = 1'b0;
wire vcc = 1'b1;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
// synopsys translate_off
initial $sdf_annotate("fir_top_v.sdo");
// synopsys translate_on

wire nx38664z1;
wire nx38664z3;
wire nx38664z9;
wire nx4119z3;
wire nx4119z2;
wire nx4119z10;
wire nx4119z12;
wire nx4119z11;
wire nx4119z9;
wire nx4119z13;
wire nx4119z15;
wire \u_audio_dac_p1_altpll|pll~clk ;
wire \u_audio_dac_p1_altpll|pll~CLK2 ;
wire audio_out_5_;
wire audio_out_4_;
wire nx24999z3;
wire audio_out_1_;
wire audio_out_0_;
wire nx24999z5;
wire audio_out_15_;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z8 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z4 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z8 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_2_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_3__dup_193 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_4__dup_192 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_6__dup_190 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_8__dup_188 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z6 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_2_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_5__dup_191 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_7__dup_189 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_8__dup_188 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|taps_16__9_ ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_17_filter_block_tap_next_7_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_9_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_5_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_3_ ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z6 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z3 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z6 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z4 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|b_10_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_9__dup_187 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z4 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_9__dup_187 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z5 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z2 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z5 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z3 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z5 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z3 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z3 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_10__dup_186 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_12_ ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z4 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_12_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z3 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_13_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z4 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z3 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z2 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z3 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z2 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z2 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z2 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z2 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z2 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_11__dup_185 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z2 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z2 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_14_ ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_12_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z2 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z2 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_ ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z2 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z4 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z1 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z17 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z9 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z13 ;
wire nx50205z4;
wire nx50205z3;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z17 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx1963z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z13 ;
wire \u_i2c_av_config|u0|nx44942z8 ;
wire \u_i2c_av_config|u0|nx7286z2 ;
wire u_sine_address_0_;
wire \u_sine_address_add9_0i1|nx37973z1 ;
wire u_sine_address_4_;
wire u_sine_address_5_;
wire u_sine_address_7_;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx51271z1 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx53265z1 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx55259z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z23 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx52268z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx55259z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx57253z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z2 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_5_ ;
wire \u_i2c_av_config|modgen_counter_cont|q_6_ ;
wire \u_i2c_av_config|nx35560z2 ;
wire \u_i2c_av_config|u0|nx22137z2 ;
wire \u_i2c_av_config|u0|sdo_5n5s2f1_0_ ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1 ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx40964z1 ;
wire \u_i2c_av_config|u0|nx41315z4 ;
wire \u_i2c_av_config|u0|nx41315z10 ;
wire \u_i2c_av_config|u0|nx41315z12 ;
wire \u_i2c_av_config|u0|nx41315z14 ;
wire \u_i2c_av_config|u0|nx41315z13 ;
wire \u_i2c_av_config|u0|nx41315z16 ;
wire \u_i2c_av_config|u0|nx41315z17 ;
wire \u_i2c_av_config|u0|nx41315z15 ;
wire \u_i2c_av_config|u0|nx41315z11 ;
wire \u_i2c_av_config|u0|nx41315z21 ;
wire \u_i2c_av_config|u0|nx41315z22 ;
wire \u_i2c_av_config|u0|nx41315z20 ;
wire \u_i2c_av_config|modgen_counter_cont|nx56256z1 ;
wire \u_i2c_av_config|modgen_counter_cont|nx57253z1 ;
wire \aud_bclk_dup0~clkctrl_outclk ;
wire \audio_out_0_~feeder_combout ;
wire \audio_out_15_~feeder_combout ;
wire nx49625z3;
wire nx49625z1;
wire nx55607z1;
wire nx49625z4;
wire display_freq_0_;
wire display_freq_1_;
wire nx49625z2;
wire display_freq_2_;
wire nx55607z2;
wire hex4_dup0_0_;
wire display_freq_3_;
wire hex4_dup0_1_;
wire hex4_dup0_2_;
wire hex4_dup0_3_;
wire hex4_dup0_4_;
wire hex4_dup0_5_;
wire hex4_dup0_6_;
wire nx38664z8;
wire display_freq_4_;
wire nx38664z2;
wire display_freq_7_;
wire nx38664z5;
wire nx38664z4;
wire display_freq_6_;
wire nx38664z6;
wire nx38664z7;
wire display_freq_5_;
wire hex5_dup0_0_;
wire hex5_dup0_1_;
wire hex5_dup0_2_;
wire hex5_dup0_3_;
wire hex5_dup0_4_;
wire hex5_dup0_5_;
wire hex5_dup0_6_;
wire nx4119z7;
wire nx4119z6;
wire nx4119z5;
wire display_freq_10_;
wire nx4119z14;
wire display_freq_8_;
wire nx4119z8;
wire display_freq_9_;
wire nx4119z1;
wire nx4119z4;
wire display_freq_11_;
wire hex6_dup0_0_;
wire hex6_dup0_1_;
wire hex6_dup0_2_;
wire hex6_dup0_3_;
wire hex6_dup0_4_;
wire hex6_dup0_5_;
wire hex6_dup0_6_;
wire nx17637z1;
wire hex7_dup0_0_;
wire \clock_27~combout ;
wire \u_audio_dac_p1_altpll|_clk1 ;
wire \u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ;
wire NOT_bit_position_0_;
wire bit_position_0_;
wire nx49817z1;
wire bit_position_2_;
wire nx48820z1;
wire bit_position_3_;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z16 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx52268z1 ;
wire nx48238z1;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z15 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z14 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z12 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx54262z1 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z11 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z10 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z8 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx56256z1 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z7 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z6 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx57253z1 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z5 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z4 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx58250z1 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z3 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z2 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z1 ;
wire \u_audio_dac_modgen_counter_lrck_1x_div|nx2038z1 ;
wire nx50205z2;
wire nx50205z1;
wire aud_adclrck_dup0;
wire \aud_adclrck_dup0~clkctrl_outclk ;
wire u_sine_address_3_;
wire \u_sine_address_add9_0i1|nx45949z23 ;
wire \u_sine_address_add9_0i1|nx38970z1 ;
wire u_sine_address_1_;
wire \u_sine_address_add9_0i1|nx45949z20 ;
wire \u_sine_address_add9_0i1|nx39967z1 ;
wire u_sine_address_2_;
wire \u_sine_address_add9_0i1|nx45949z17 ;
wire \u_sine_address_add9_0i1|nx40964z1 ;
wire \u_sine_address_add9_0i1|nx45949z14 ;
wire \u_sine_address_add9_0i1|nx41961z1 ;
wire \u_sine_address_add9_0i1|nx45949z11 ;
wire \u_sine_address_add9_0i1|nx42958z1 ;
wire u_sine_address_6_;
wire \u_sine_address_add9_0i1|nx45949z8 ;
wire \u_sine_address_add9_0i1|nx43955z1 ;
wire \u_sine_address_add9_0i1|nx45949z5 ;
wire \u_sine_address_add9_0i1|nx44952z1 ;
wire u_sine_address_8_;
wire \u_sine_address_add9_0i1|nx45949z3 ;
wire \u_sine_address_add9_0i1|nx45949z1 ;
wire \u_noise_modgen_counter_address|nx51271z1 ;
wire \u_noise_modgen_counter_address|q_0_ ;
wire \u_noise_modgen_counter_address|nx60244z10 ;
wire \u_noise_modgen_counter_address|nx52268z1 ;
wire \u_noise_modgen_counter_address|q_1_ ;
wire \u_noise_modgen_counter_address|nx60244z9 ;
wire \u_noise_modgen_counter_address|nx53265z1 ;
wire \u_noise_modgen_counter_address|q_2_ ;
wire \u_noise_modgen_counter_address|nx60244z8 ;
wire \u_noise_modgen_counter_address|nx54262z1 ;
wire \u_noise_modgen_counter_address|q_3_ ;
wire \u_noise_modgen_counter_address|nx60244z7 ;
wire \u_noise_modgen_counter_address|nx55259z1 ;
wire \u_noise_modgen_counter_address|q_4_ ;
wire \u_noise_modgen_counter_address|nx60244z6 ;
wire \u_noise_modgen_counter_address|nx56256z1 ;
wire \u_noise_modgen_counter_address|q_5_ ;
wire \u_noise_modgen_counter_address|nx60244z5 ;
wire \u_noise_modgen_counter_address|nx57253z1 ;
wire \u_noise_modgen_counter_address|q_6_ ;
wire \u_noise_modgen_counter_address|nx60244z4 ;
wire \u_noise_modgen_counter_address|nx58250z1 ;
wire \u_noise_modgen_counter_address|q_7_ ;
wire \u_noise_modgen_counter_address|nx60244z3 ;
wire \u_noise_modgen_counter_address|nx59247z1 ;
wire \u_noise_modgen_counter_address|q_8_ ;
wire \u_noise_modgen_counter_address|nx60244z2 ;
wire \u_noise_modgen_counter_address|nx60244z1 ;
wire \u_noise_modgen_counter_address|q_9_ ;
wire raw_audio_9_;
wire raw_audio_11_;
wire \u_fir|taps_1__15_ ;
wire \u_fir|taps_2__15_ ;
wire \u_fir|taps_3__15_ ;
wire \u_fir|taps_4__15_ ;
wire \u_fir|taps_5__15_ ;
wire \u_fir|taps_6__15_ ;
wire \u_fir|taps_7__15_ ;
wire \u_fir|taps_8__15_ ;
wire \u_fir|taps_9__15_ ;
wire \u_fir|taps_10__15_ ;
wire \u_fir|taps_11__15_ ;
wire \u_fir|taps_12__15_ ;
wire raw_audio_10_;
wire \u_fir|taps_1__10_ ;
wire \u_fir|taps_2__10_ ;
wire \u_fir|taps_3__10_~feeder_combout ;
wire \u_fir|taps_3__10_ ;
wire \u_fir|taps_4__10_ ;
wire \u_fir|taps_5__10_ ;
wire \u_fir|taps_6__10_ ;
wire \u_fir|taps_7__10_ ;
wire \u_fir|taps_8__10_ ;
wire \u_fir|taps_9__10_ ;
wire \u_fir|taps_10__10_ ;
wire \u_fir|taps_11__10_ ;
wire \u_fir|taps_12__10_ ;
wire raw_audio_8_;
wire \u_fir|taps_1__8_ ;
wire \u_fir|taps_2__8_ ;
wire \u_fir|taps_3__8_~feeder_combout ;
wire \u_fir|taps_3__8_ ;
wire \u_fir|taps_4__8_ ;
wire \u_fir|taps_5__8_ ;
wire \u_fir|taps_6__8_ ;
wire \u_fir|taps_7__8_ ;
wire \u_fir|taps_8__8_ ;
wire \u_fir|taps_9__8_ ;
wire \u_fir|taps_10__8_ ;
wire \u_fir|taps_11__8_ ;
wire \u_fir|taps_12__8_ ;
wire raw_audio_7_;
wire \u_fir|taps_1__7_ ;
wire \u_fir|taps_2__7_ ;
wire \u_fir|taps_3__7_~feeder_combout ;
wire \u_fir|taps_3__7_ ;
wire \u_fir|taps_4__7_ ;
wire \u_fir|taps_5__7_ ;
wire \u_fir|taps_6__7_ ;
wire \u_fir|taps_7__7_ ;
wire \u_fir|taps_8__7_ ;
wire \u_fir|taps_9__7_ ;
wire \u_fir|taps_10__7_ ;
wire \u_fir|taps_11__7_ ;
wire \u_fir|taps_12__7_ ;
wire raw_audio_5_;
wire \u_fir|taps_1__5_ ;
wire \u_fir|taps_2__5_ ;
wire \u_fir|taps_3__5_~feeder_combout ;
wire \u_fir|taps_3__5_ ;
wire \u_fir|taps_4__5_ ;
wire \u_fir|taps_5__5_ ;
wire \u_fir|taps_6__5_ ;
wire \u_fir|taps_7__5_ ;
wire \u_fir|taps_8__5_ ;
wire \u_fir|taps_9__5_ ;
wire \u_fir|taps_10__5_ ;
wire \u_fir|taps_11__5_ ;
wire \u_fir|taps_12__5_ ;
wire raw_audio_3_;
wire \u_fir|taps_1__3_~feeder_combout ;
wire \u_fir|taps_1__3_ ;
wire \u_fir|taps_2__3_ ;
wire \u_fir|taps_3__3_ ;
wire \u_fir|taps_4__3_ ;
wire \u_fir|taps_5__3_ ;
wire \u_fir|taps_6__3_~feeder_combout ;
wire \u_fir|taps_6__3_ ;
wire \u_fir|taps_7__3_~feeder_combout ;
wire \u_fir|taps_7__3_ ;
wire \u_fir|taps_8__3_ ;
wire \u_fir|taps_9__3_ ;
wire \u_fir|taps_10__3_ ;
wire \u_fir|taps_11__3_ ;
wire \u_fir|taps_12__3_ ;
wire raw_audio_1_;
wire \u_fir|taps_1__1_ ;
wire \u_fir|taps_2__1_ ;
wire \u_fir|taps_3__1_ ;
wire \u_fir|taps_4__1_ ;
wire \u_fir|taps_5__1_~feeder_combout ;
wire \u_fir|taps_5__1_ ;
wire \u_fir|taps_6__1_~feeder_combout ;
wire \u_fir|taps_6__1_ ;
wire \u_fir|taps_7__1_~feeder_combout ;
wire \u_fir|taps_7__1_ ;
wire \u_fir|taps_8__1_ ;
wire \u_fir|taps_9__1_ ;
wire \u_fir|taps_10__1_ ;
wire \u_fir|taps_11__1_ ;
wire \u_fir|taps_12__1_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z16 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z15 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z13 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z11 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z9 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z7 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z6 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|b_10_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z5 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_ ;
wire raw_audio_6_;
wire \u_fir|taps_1__6_ ;
wire \u_fir|taps_2__6_ ;
wire \u_fir|taps_3__6_~feeder_combout ;
wire \u_fir|taps_3__6_ ;
wire \u_fir|taps_4__6_ ;
wire \u_fir|taps_5__6_ ;
wire \u_fir|taps_6__6_ ;
wire \u_fir|taps_7__6_ ;
wire \u_fir|taps_8__6_ ;
wire \u_fir|taps_9__6_ ;
wire \u_fir|taps_10__6_ ;
wire \u_fir|taps_11__6_ ;
wire \u_fir|taps_12__6_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_4_ ;
wire raw_audio_0_;
wire \u_fir|taps_1__0_ ;
wire \u_fir|taps_2__0_~feeder_combout ;
wire \u_fir|taps_2__0_ ;
wire \u_fir|taps_3__0_~feeder_combout ;
wire \u_fir|taps_3__0_ ;
wire \u_fir|taps_4__0_ ;
wire \u_fir|taps_5__0_ ;
wire \u_fir|taps_6__0_~feeder_combout ;
wire \u_fir|taps_6__0_ ;
wire \u_fir|taps_7__0_ ;
wire \u_fir|taps_8__0_ ;
wire \u_fir|taps_9__0_ ;
wire \u_fir|taps_10__0_~feeder_combout ;
wire \u_fir|taps_10__0_ ;
wire \u_fir|taps_11__0_~feeder_combout ;
wire \u_fir|taps_11__0_ ;
wire \u_fir|taps_12__0_ ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z26 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z25 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z23 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z21 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z19 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z17 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z4 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z3 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_ ;
wire \u_fir|taps_1__9_ ;
wire \u_fir|taps_2__9_ ;
wire \u_fir|taps_3__9_~feeder_combout ;
wire \u_fir|taps_3__9_ ;
wire \u_fir|taps_4__9_ ;
wire \u_fir|taps_5__9_ ;
wire \u_fir|taps_6__9_ ;
wire \u_fir|taps_7__9_ ;
wire \u_fir|taps_8__9_ ;
wire \u_fir|taps_9__9_ ;
wire \u_fir|taps_10__9_ ;
wire \u_fir|taps_11__9_ ;
wire raw_audio_4_;
wire \u_fir|taps_1__4_ ;
wire \u_fir|taps_2__4_ ;
wire \u_fir|taps_3__4_ ;
wire \u_fir|taps_4__4_ ;
wire \u_fir|taps_5__4_ ;
wire \u_fir|taps_6__4_ ;
wire \u_fir|taps_7__4_ ;
wire \u_fir|taps_8__4_ ;
wire \u_fir|taps_9__4_ ;
wire \u_fir|taps_10__4_ ;
wire \u_fir|taps_11__4_ ;
wire raw_audio_2_;
wire \u_fir|taps_1__2_ ;
wire \u_fir|taps_2__2_ ;
wire \u_fir|taps_3__2_ ;
wire \u_fir|taps_4__2_ ;
wire \u_fir|taps_5__2_~feeder_combout ;
wire \u_fir|taps_5__2_ ;
wire \u_fir|taps_6__2_~feeder_combout ;
wire \u_fir|taps_6__2_ ;
wire \u_fir|taps_7__2_~feeder_combout ;
wire \u_fir|taps_7__2_ ;
wire \u_fir|taps_8__2_ ;
wire \u_fir|taps_9__2_ ;
wire \u_fir|taps_10__2_ ;
wire \u_fir|taps_11__2_ ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z13 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z12 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z10 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z8 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z6 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z4 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z3 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z13 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z12 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z10 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z8 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z13 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z12 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z10 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z8 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z16 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z15 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z13 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z11 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z26 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z25 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z23 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_5__dup_191 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z13 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z12 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z10 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z13 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z12 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z10 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_11_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192 ;
wire \u_fir|tap_array_12_filter_block_prod_mults28_0|d_3__dup_193 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|taps_13__15_ ;
wire \u_fir|taps_12__9_ ;
wire \u_fir|taps_13__9_ ;
wire \u_fir|taps_13__8_ ;
wire \u_fir|taps_13__7_ ;
wire \u_fir|taps_12__4_ ;
wire \u_fir|taps_13__4_ ;
wire \u_fir|taps_13__5_ ;
wire \u_fir|taps_12__2_ ;
wire \u_fir|taps_13__2_ ;
wire \u_fir|taps_13__1_ ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z13 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z12 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z10 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z8 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z6 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z4 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z3 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_13_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|taps_13__10_ ;
wire \u_fir|taps_14__10_ ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|taps_14__7_ ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|taps_14__5_ ;
wire \u_fir|taps_14__4_ ;
wire \u_fir|taps_13__3_ ;
wire \u_fir|taps_14__3_ ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|taps_14__15_ ;
wire \u_fir|taps_15__15_ ;
wire \u_fir|taps_14__9_ ;
wire \u_fir|taps_15__9_ ;
wire \u_fir|taps_15__7_ ;
wire \u_fir|taps_14__8_ ;
wire \u_fir|taps_15__8_ ;
wire \u_fir|taps_15__4_ ;
wire \u_fir|taps_13__6_ ;
wire \u_fir|taps_14__6_ ;
wire \u_fir|taps_15__6_ ;
wire \u_fir|taps_14__2_ ;
wire \u_fir|taps_15__2_ ;
wire \u_fir|taps_14__1_~feeder_combout ;
wire \u_fir|taps_14__1_ ;
wire \u_fir|taps_15__1_ ;
wire \u_fir|taps_15__3_ ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z17 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z16 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z15 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z14 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z12 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z10 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z8 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z6 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z5 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_13_ ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx41961z1 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx37973z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|taps_15__10_ ;
wire \u_fir|taps_16__10_ ;
wire \u_fir|taps_16__8_ ;
wire \u_fir|taps_16__7_ ;
wire \u_fir|taps_15__5_ ;
wire \u_fir|taps_16__5_ ;
wire \u_fir|taps_16__3_ ;
wire \u_fir|taps_16__1_ ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z13 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z12 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z11 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z10 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z8 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z6 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z4 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z3 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z2 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_16_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_17_filter_block_tap_next_10_ ;
wire \u_fir|taps_16__15_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_15_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_8_ ;
wire \u_fir|taps_16__6_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_6_ ;
wire \u_fir|taps_16__4_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_4_ ;
wire \u_fir|taps_16__2_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_2_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_1_ ;
wire \u_fir|taps_13__0_ ;
wire \u_fir|taps_14__0_~feeder_combout ;
wire \u_fir|taps_14__0_ ;
wire \u_fir|taps_15__0_ ;
wire \u_fir|taps_16__0_ ;
wire \u_fir|tap_array_17_filter_block_tap_next_0_ ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z15 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z14 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z12 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z10 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z8 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z6 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z5 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx46946z1 ;
wire audio_out_9_;
wire nx50814z1;
wire bit_position_1_;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx45949z1 ;
wire audio_out_8_;
wire nx24999z7;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z4 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z3 ;
wire \u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_ ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx62798z1 ;
wire audio_out_10_;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx63795z1 ;
wire audio_out_11_;
wire nx24999z6;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx44952z1 ;
wire audio_out_7_;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx43955z1 ;
wire audio_out_6_;
wire nx24999z2;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx40964z1 ;
wire audio_out_3_;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx39967z1 ;
wire audio_out_2_;
wire nx24999z4;
wire nx24999z1;
wire \audio_out_13_~feeder_combout ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z4 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z3 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z2 ;
wire \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z6 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z4 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z3 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z2 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z9 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z7 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z6 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z21 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z19 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z17 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z4 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_11__dup_185 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z13 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z12 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z10 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z8 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z6 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z13 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z12 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z11 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z10 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z8 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z6 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5 ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_2_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z15 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z14 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z12 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z10 ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_ ;
wire \u_fir|tap_array_1_filter_block_prod_mults28_0|d_3_ ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z17 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z16 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z15 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z14 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z12 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z10 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_3_filter_block_prod_mults28_0|d_5_ ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_ ;
wire \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx39967z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z43 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_6_filter_block_prod_mults28_0|d_7__dup_189 ;
wire \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7 ;
wire \u_fir|tap_array_7_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z8 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z6 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z4 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_ ;
wire \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx43955z1 ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_ ;
wire \u_fir|tap_array_8_filter_block_prod_mults28_0|d_7_ ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z37 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx45949z1 ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_9_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z8 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z6 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z4 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z3 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_11_ ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1 ;
wire \u_fir|tap_array_10_filter_block_prod_mults28_0|d_9_ ;
wire \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z31 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z25 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx62798z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z19 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx64792z1 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z13 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx253z1 ;
wire audio_out_13_;
wire \audio_out_12_~feeder_combout ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx64792z1 ;
wire audio_out_12_;
wire nx24999z9;
wire \audio_out_14_~feeder_combout ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx1250z1 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z7 ;
wire \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx1250z1 ;
wire audio_out_14_;
wire nx24999z8;
wire aud_dacdat_dup0;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z10 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx52268z1 ;
wire \u_i2c_av_config|modgen_counter_cont|nx51271z1 ;
wire \u_i2c_av_config|modgen_counter_cont|nx17096z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_10_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx59247z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_8_ ;
wire \u_i2c_av_config|nx35560z3 ;
wire \u_i2c_av_config|modgen_counter_cont|nx54262z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_3_ ;
wire \u_i2c_av_config|nx17807z2 ;
wire \u_i2c_av_config|nx35560z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_0_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z16 ;
wire \u_i2c_av_config|modgen_counter_cont|nx52268z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_1_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z15 ;
wire \u_i2c_av_config|modgen_counter_cont|nx53265z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_2_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z14 ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z13 ;
wire \u_i2c_av_config|modgen_counter_cont|nx55259z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_4_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z12 ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z11 ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z10 ;
wire \u_i2c_av_config|modgen_counter_cont|nx58250z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_7_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z9 ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z8 ;
wire \u_i2c_av_config|modgen_counter_cont|nx60244z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_9_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z7 ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z6 ;
wire \u_i2c_av_config|modgen_counter_cont|nx18093z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_11_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z5 ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z4 ;
wire \u_i2c_av_config|modgen_counter_cont|nx20087z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_13_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z3 ;
wire \u_i2c_av_config|modgen_counter_cont|nx21084z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_14_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z2 ;
wire \u_i2c_av_config|modgen_counter_cont|nx22081z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_15_ ;
wire \u_i2c_av_config|modgen_counter_cont|nx19090z1 ;
wire \u_i2c_av_config|modgen_counter_cont|q_12_ ;
wire \u_i2c_av_config|nx35560z4 ;
wire \u_i2c_av_config|nx17807z1 ;
wire \u_i2c_av_config|reset_n ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx51271z1 ;
wire \u_i2c_av_config|nx23875z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z25 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z24 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z22 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx53265z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z21 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z20 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z18 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z16 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx56256z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z15 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z14 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z12 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx58250z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z11 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z10 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx59247z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z9 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z8 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx60244z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z7 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z6 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z4 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx18093z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3 ;
wire \u_i2c_av_config|nx2692z4 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx54262z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z19 ;
wire \u_i2c_av_config|nx2692z3 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx17096z1 ;
wire \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z5 ;
wire \u_i2c_av_config|nx2692z5 ;
wire \u_i2c_av_config|nx2692z2 ;
wire \u_i2c_av_config|nx2692z1 ;
wire \u_i2c_av_config|m_i2c_ctrl_clk ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z2 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z1 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx51271z1 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ;
wire \u_i2c_av_config|u0|nx7286z1 ;
wire \u_i2c_av_config|nx51161z1 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z8 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z6 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx54262z1 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z4 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z1 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx53265z1 ;
wire \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ;
wire \u_i2c_av_config|u0|nx43379z2 ;
wire \u_i2c_av_config|u0|nx43379z4 ;
wire \u_i2c_av_config|u0|nx43379z3 ;
wire \u_i2c_av_config|u0|nx44942z1 ;
wire \u_i2c_av_config|u0|nx44942z7 ;
wire \u_i2c_av_config|u0|nx44942z6 ;
wire \u_i2c_av_config|u0|nx44942z5 ;
wire \u_i2c_av_config|u0|nx44942z3 ;
wire \u_i2c_av_config|u0|nx44942z2 ;
wire \u_i2c_av_config|u0|nx43379z1 ;
wire \u_i2c_av_config|u0|p_i2c_sclk ;
wire \clock_27~clkctrl_outclk ;
wire \u_i2c_av_config|u0|sdo_5n5s2f1_1_ ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11 ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z8 ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z5 ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z3 ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1 ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1 ;
wire \u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1 ;
wire \u_i2c_av_config|u0|nx41315z18 ;
wire \u_i2c_av_config|u0|nx41315z9 ;
wire \u_i2c_av_config|u0|nx44942z4 ;
wire \u_i2c_av_config|u0|nx41315z5 ;
wire \u_i2c_av_config|u0|nx41315z6 ;
wire \u_i2c_av_config|u0|nx22137z1 ;
wire \u_i2c_av_config|u0|nx41315z3 ;
wire \u_i2c_av_config|u0|nx41315z8 ;
wire \u_i2c_av_config|u0|nx41315z2 ;
wire \u_i2c_av_config|u0|nx41315z7 ;
wire \u_i2c_av_config|u0|nx41315z1 ;
wire \u_i2c_av_config|u0|nx41315z19 ;
wire \u_i2c_av_config|u0|nx51857z1 ;
wire nx30102z1;
wire nx30102z2;
wire u_audio_dac_bck_div_2_;
wire nx32096z1;
wire u_audio_dac_bck_div_0_;
wire nx31099z1;
wire nx31099z2;
wire u_audio_dac_bck_div_1_;
wire nx15494z1;
wire aud_bclk_dup0;
wire [11:0] \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a ;
wire [7:0] \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a ;
wire [3:0] \key~combout ;
wire [17:0] \sw~combout ;

wire [2:0] \u_audio_dac_p1_altpll|pll_CLK_bus ;
wire [3:0] \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0_PORTADATAOUT_bus ;
wire [11:0] \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus ;
wire [3:0] \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4_PORTADATAOUT_bus ;

assign \u_audio_dac_p1_altpll|pll~clk  = \u_audio_dac_p1_altpll|pll_CLK_bus [0];
assign \u_audio_dac_p1_altpll|_clk1  = \u_audio_dac_p1_altpll|pll_CLK_bus [1];
assign \u_audio_dac_p1_altpll|pll~CLK2  = \u_audio_dac_p1_altpll|pll_CLK_bus [2];

assign \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [0] = \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0_PORTADATAOUT_bus [0];
assign \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [1] = \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0_PORTADATAOUT_bus [1];
assign \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [2] = \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0_PORTADATAOUT_bus [2];
assign \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [3] = \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0_PORTADATAOUT_bus [3];

assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [0] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [0];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [1] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [1];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [2] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [2];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [3] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [3];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [4] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [4];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [5] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [5];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [6] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [6];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [7] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [7];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [8] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [8];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [9] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [9];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [10] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [10];
assign \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [11] = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus [11];

assign \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [4] = \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4_PORTADATAOUT_bus [0];
assign \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [5] = \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4_PORTADATAOUT_bus [1];
assign \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [6] = \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4_PORTADATAOUT_bus [2];
assign \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [7] = \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4_PORTADATAOUT_bus [3];

// atom is at LCCOMB_X31_Y14_N10
cycloneii_lcell_comb ix38664z52925(
// Equation(s):
// nx38664z1 = \sw~combout [3] & (!\sw~combout [1] & \sw~combout [4]) # !\sw~combout [3] & \sw~combout [0] & \sw~combout [1] & !\sw~combout [4]

	.dataa(\sw~combout [3]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [1]),
	.datad(\sw~combout [4]),
	.cin(gnd),
	.combout(nx38664z1),
	.cout());
// synopsys translate_off
defparam ix38664z52925.lut_mask = 16'h0A40;
defparam ix38664z52925.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N16
cycloneii_lcell_comb ix38664z52928(
// Equation(s):
// nx38664z3 = \sw~combout [1] & (\sw~combout [2] $ (\sw~combout [0] & !\sw~combout [3])) # !\sw~combout [1] & \sw~combout [2] & (\sw~combout [0] # !\sw~combout [3])

	.dataa(\sw~combout [1]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx38664z3),
	.cout());
// synopsys translate_off
defparam ix38664z52928.lut_mask = 16'hE708;
defparam ix38664z52928.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N2
cycloneii_lcell_comb ix38664z52936(
// Equation(s):
// nx38664z9 = \sw~combout [4] & !\sw~combout [2] & (\sw~combout [5] # !\sw~combout [6]) # !\sw~combout [4] & (\sw~combout [2])

	.dataa(\sw~combout [5]),
	.datab(\sw~combout [6]),
	.datac(\sw~combout [4]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx38664z9),
	.cout());
// synopsys translate_off
defparam ix38664z52936.lut_mask = 16'h0FB0;
defparam ix38664z52936.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N8
cycloneii_lcell_comb ix4119z52927(
// Equation(s):
// nx4119z3 = !\sw~combout [2] & !\sw~combout [0] & !\sw~combout [4] & !\sw~combout [1]

	.dataa(\sw~combout [2]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [4]),
	.datad(\sw~combout [1]),
	.cin(gnd),
	.combout(nx4119z3),
	.cout());
// synopsys translate_off
defparam ix4119z52927.lut_mask = 16'h0001;
defparam ix4119z52927.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N10
cycloneii_lcell_comb ix4119z52926(
// Equation(s):
// nx4119z2 = \sw~combout [5] & (nx4119z3) # !\sw~combout [5] & \sw~combout [4]

	.dataa(vcc),
	.datab(\sw~combout [4]),
	.datac(\sw~combout [5]),
	.datad(nx4119z3),
	.cin(gnd),
	.combout(nx4119z2),
	.cout());
// synopsys translate_off
defparam ix4119z52926.lut_mask = 16'hFC0C;
defparam ix4119z52926.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N0
cycloneii_lcell_comb ix4119z52936(
// Equation(s):
// nx4119z10 = \sw~combout [5] & (\sw~combout [1] & \sw~combout [2]) # !\sw~combout [5] & !\sw~combout [6]

	.dataa(\sw~combout [5]),
	.datab(\sw~combout [6]),
	.datac(\sw~combout [1]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx4119z10),
	.cout());
// synopsys translate_off
defparam ix4119z52936.lut_mask = 16'hB111;
defparam ix4119z52936.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N26
cycloneii_lcell_comb ix4119z52938(
// Equation(s):
// nx4119z12 = \sw~combout [5] & !\sw~combout [0] & !\sw~combout [1] & !\sw~combout [2]

	.dataa(\sw~combout [5]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [1]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx4119z12),
	.cout());
// synopsys translate_off
defparam ix4119z52938.lut_mask = 16'h0002;
defparam ix4119z52938.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N4
cycloneii_lcell_comb ix4119z52937(
// Equation(s):
// nx4119z11 = \sw~combout [4] # \sw~combout [6] & !\sw~combout [5] # !\sw~combout [6] & (nx4119z12)

	.dataa(\sw~combout [5]),
	.datab(\sw~combout [4]),
	.datac(\sw~combout [6]),
	.datad(nx4119z12),
	.cin(gnd),
	.combout(nx4119z11),
	.cout());
// synopsys translate_off
defparam ix4119z52937.lut_mask = 16'hDFDC;
defparam ix4119z52937.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N30
cycloneii_lcell_comb ix4119z52935(
// Equation(s):
// nx4119z9 = nx4119z11 & (nx4119z10 # !\sw~combout [4])

	.dataa(vcc),
	.datab(nx4119z11),
	.datac(\sw~combout [4]),
	.datad(nx4119z10),
	.cin(gnd),
	.combout(nx4119z9),
	.cout());
// synopsys translate_off
defparam ix4119z52935.lut_mask = 16'hCC0C;
defparam ix4119z52935.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N6
cycloneii_lcell_comb ix4119z52940(
// Equation(s):
// nx4119z13 = \sw~combout [5] $ (\sw~combout [2] & \sw~combout [3] & \sw~combout [1] # !\sw~combout [2] & !\sw~combout [3])

	.dataa(\sw~combout [2]),
	.datab(\sw~combout [5]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [1]),
	.cin(gnd),
	.combout(nx4119z13),
	.cout());
// synopsys translate_off
defparam ix4119z52940.lut_mask = 16'h69C9;
defparam ix4119z52940.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N24
cycloneii_lcell_comb ix4119z52942(
// Equation(s):
// nx4119z15 = \sw~combout [5] $ (\sw~combout [2] # \sw~combout [0] # \sw~combout [1])

	.dataa(\sw~combout [2]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [5]),
	.datad(\sw~combout [1]),
	.cin(gnd),
	.combout(nx4119z15),
	.cout());
// synopsys translate_off
defparam ix4119z52942.lut_mask = 16'h0F1E;
defparam ix4119z52942.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y14_N1
cycloneii_lcell_ff reg_audio_out_5_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_5_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx42958z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_5_));

// atom is at LCFF_X34_Y14_N3
cycloneii_lcell_ff reg_audio_out_4_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_4_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx41961z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_4_));

// atom is at LCCOMB_X34_Y14_N14
cycloneii_lcell_comb ix24999z52926(
// Equation(s):
// nx24999z3 = bit_position_0_ & (bit_position_1_ & audio_out_4_) # !bit_position_0_ & (audio_out_5_ # !bit_position_1_)

	.dataa(bit_position_0_),
	.datab(audio_out_5_),
	.datac(bit_position_1_),
	.datad(audio_out_4_),
	.cin(gnd),
	.combout(nx24999z3),
	.cout());
// synopsys translate_off
defparam ix24999z52926.lut_mask = 16'hE545;
defparam ix24999z52926.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y14_N5
cycloneii_lcell_ff reg_audio_out_1_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_1_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx38970z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_1_));

// atom is at LCFF_X34_Y14_N7
cycloneii_lcell_ff reg_audio_out_0_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\audio_out_0_~feeder_combout ),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx37973z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_0_));

// atom is at LCCOMB_X34_Y14_N8
cycloneii_lcell_comb ix24999z52928(
// Equation(s):
// nx24999z5 = bit_position_1_ & (bit_position_0_ & audio_out_0_ # !bit_position_0_ & (audio_out_1_)) # !bit_position_1_ & (!bit_position_0_)

	.dataa(audio_out_0_),
	.datab(bit_position_1_),
	.datac(audio_out_1_),
	.datad(bit_position_0_),
	.cin(gnd),
	.combout(nx24999z5),
	.cout());
// synopsys translate_off
defparam ix24999z52928.lut_mask = 16'h88F3;
defparam ix24999z52928.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X35_Y14_N11
cycloneii_lcell_ff reg_audio_out_15_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\audio_out_15_~feeder_combout ),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_15_));

// atom is at LCCOMB_X48_Y16_N12
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52932 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_1__6_  $ \u_fir|taps_1__9_  $ !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z10 ) # GND
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9  = CARRY(\u_fir|taps_1__6_  & (\u_fir|taps_1__9_  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z10 ) # !\u_fir|taps_1__6_  & \u_fir|taps_1__9_  & 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z10 )

	.dataa(\u_fir|taps_1__6_ ),
	.datab(\u_fir|taps_1__9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z10 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N14
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52931 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_1__10_  & (\u_fir|taps_1__7_  & \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9  & VCC # !\u_fir|taps_1__7_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9 ) # 
// !\u_fir|taps_1__10_  & (\u_fir|taps_1__7_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9  # !\u_fir|taps_1__7_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9  # GND))
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z8  = CARRY(\u_fir|taps_1__10_  & !\u_fir|taps_1__7_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9  # !\u_fir|taps_1__10_  & (!\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9  # 
// !\u_fir|taps_1__7_ ))

	.dataa(\u_fir|taps_1__10_ ),
	.datab(\u_fir|taps_1__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z9 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N16
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52930 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_1__8_  $ \u_fir|taps_1__15_  $ !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z8 ) # GND
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7  = CARRY(\u_fir|taps_1__8_  & (\u_fir|taps_1__15_  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z8 ) # !\u_fir|taps_1__8_  & \u_fir|taps_1__15_  & 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z8 )

	.dataa(\u_fir|taps_1__8_ ),
	.datab(\u_fir|taps_1__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z8 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N8
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52932 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_2__4_  $ \u_fir|taps_2__5_  $ !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z10 ) # GND
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9  = CARRY(\u_fir|taps_2__4_  & (\u_fir|taps_2__5_  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z10 ) # !\u_fir|taps_2__4_  & \u_fir|taps_2__5_  & 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z10 )

	.dataa(\u_fir|taps_2__4_ ),
	.datab(\u_fir|taps_2__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z10 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N10
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52931 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_2__6_  & (\u_fir|taps_2__5_  & \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9  & VCC # !\u_fir|taps_2__5_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9 ) # 
// !\u_fir|taps_2__6_  & (\u_fir|taps_2__5_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9  # !\u_fir|taps_2__5_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9  # GND))
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z8  = CARRY(\u_fir|taps_2__6_  & !\u_fir|taps_2__5_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9  # !\u_fir|taps_2__6_  & (!\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9  # 
// !\u_fir|taps_2__5_ ))

	.dataa(\u_fir|taps_2__6_ ),
	.datab(\u_fir|taps_2__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z9 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N12
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52930 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_2__7_  $ \u_fir|taps_2__6_  $ !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z8 ) # GND
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7  = CARRY(\u_fir|taps_2__7_  & (\u_fir|taps_2__6_  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z8 ) # !\u_fir|taps_2__7_  & \u_fir|taps_2__6_  & 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z8 )

	.dataa(\u_fir|taps_2__7_ ),
	.datab(\u_fir|taps_2__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z8 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N14
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52929 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_2__7_  & (\u_fir|taps_2__8_  & \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7  & VCC # !\u_fir|taps_2__8_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7 ) # 
// !\u_fir|taps_2__7_  & (\u_fir|taps_2__8_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7  # !\u_fir|taps_2__8_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7  # GND))
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z6  = CARRY(\u_fir|taps_2__7_  & !\u_fir|taps_2__8_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7  # !\u_fir|taps_2__7_  & (!\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7  # 
// !\u_fir|taps_2__8_ ))

	.dataa(\u_fir|taps_2__7_ ),
	.datab(\u_fir|taps_2__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z7 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N18
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52927 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_2__9_  & (\u_fir|taps_2__10_  & \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5  & VCC # !\u_fir|taps_2__10_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5 ) # 
// !\u_fir|taps_2__9_  & (\u_fir|taps_2__10_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5  # !\u_fir|taps_2__10_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5  # GND))
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z4  = CARRY(\u_fir|taps_2__9_  & !\u_fir|taps_2__10_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5  # !\u_fir|taps_2__9_  & (!\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5  # 
// !\u_fir|taps_2__10_ ))

	.dataa(\u_fir|taps_2__9_ ),
	.datab(\u_fir|taps_2__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N0
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_2_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_3_  $ VCC) # !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_4_  & 
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_3_  & VCC
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_4_  & \u_fir|tap_array_1_filter_block_prod_mults28_0|d_3_ )

	.dataa(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_4_ ),
	.datab(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N2
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_2_filter_block_prod_mults28_0|d_5_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_5_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_  & 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_5_  & (!\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_ ))

	.dataa(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_5_ ),
	.datab(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N6
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_2_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_  & 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_7_  & (!\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_ ))

	.dataa(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N8
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_7_  $ \u_fir|tap_array_2_filter_block_prod_mults28_0|d_8_  $ !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|d_8_  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_7_  & \u_fir|tap_array_2_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N10
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_1_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_  & 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_8_  & (!\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_ ))

	.dataa(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_8_ ),
	.datab(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y16_N30
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52933 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_3__8_  & (\u_fir|taps_3__5_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11  # !\u_fir|taps_3__5_  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11  # GND)) # 
// !\u_fir|taps_3__8_  & (\u_fir|taps_3__5_  & \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11  & VCC # !\u_fir|taps_3__5_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11 )
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z10  = CARRY(\u_fir|taps_3__8_  & (!\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11  # !\u_fir|taps_3__5_ ) # !\u_fir|taps_3__8_  & !\u_fir|taps_3__5_  & 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11 )

	.dataa(\u_fir|taps_3__8_ ),
	.datab(\u_fir|taps_3__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52933 .lut_mask = 16'h692B;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N2
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52931 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_3__7_  & (\u_fir|taps_3__10_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9  # !\u_fir|taps_3__10_  & \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9  & VCC) # 
// !\u_fir|taps_3__7_  & (\u_fir|taps_3__10_  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9  # GND) # !\u_fir|taps_3__10_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9 )
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z8  = CARRY(\u_fir|taps_3__7_  & \u_fir|taps_3__10_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9  # !\u_fir|taps_3__7_  & (\u_fir|taps_3__10_  # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9 ))

	.dataa(\u_fir|taps_3__7_ ),
	.datab(\u_fir|taps_3__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52931 .lut_mask = 16'h694D;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N4
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52930 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_3__8_  $ \u_fir|taps_3__15_  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z8 ) # GND
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7  = CARRY(\u_fir|taps_3__8_  & (!\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z8  # !\u_fir|taps_3__15_ ) # !\u_fir|taps_3__8_  & !\u_fir|taps_3__15_  & 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z8 )

	.dataa(\u_fir|taps_3__8_ ),
	.datab(\u_fir|taps_3__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z8 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52930 .lut_mask = 16'h962B;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N0
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_5_  $ VCC) # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx37973z1  & 
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_5_  & VCC
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|tap_array_3_filter_block_prod_mults28_0|d_5_ )

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N2
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_  & \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_  & 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_ ))

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N4
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_7_  $ \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx39967z1  $ !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx39967z1  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_7_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx39967z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx39967z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N8
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|d_9_  $ !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_9_  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|tap_array_3_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N10
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_3_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_10_  & (!\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N6
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|taps_4__6_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|taps_4__6_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1  & 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|taps_4__6_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|taps_4__6_  & 
// (!\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1 ))

	.dataa(\u_fir|taps_4__6_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N8
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|taps_4__7_  $ !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|taps_4__7_  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|taps_4__7_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|taps_4__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N10
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|taps_4__8_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|taps_4__8_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|taps_4__8_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|taps_4__8_  & 
// (!\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|taps_4__8_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N10
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52933 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_5__5_  & (\u_fir|taps_5__3_  & \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11  & VCC # !\u_fir|taps_5__3_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11 ) # 
// !\u_fir|taps_5__5_  & (\u_fir|taps_5__3_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_5__3_  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11  # GND))
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z10  = CARRY(\u_fir|taps_5__5_  & !\u_fir|taps_5__3_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_5__5_  & (!\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11  # 
// !\u_fir|taps_5__3_ ))

	.dataa(\u_fir|taps_5__5_ ),
	.datab(\u_fir|taps_5__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N12
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52932 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_5__6_  $ \u_fir|taps_5__4_  $ !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z10 ) # GND
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9  = CARRY(\u_fir|taps_5__6_  & (\u_fir|taps_5__4_  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z10 ) # !\u_fir|taps_5__6_  & \u_fir|taps_5__4_  & 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z10 )

	.dataa(\u_fir|taps_5__6_ ),
	.datab(\u_fir|taps_5__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z10 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N14
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52931 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_5__5_  & (\u_fir|taps_5__7_  & \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9  & VCC # !\u_fir|taps_5__7_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9 ) # 
// !\u_fir|taps_5__5_  & (\u_fir|taps_5__7_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_5__7_  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9  # GND))
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z8  = CARRY(\u_fir|taps_5__5_  & !\u_fir|taps_5__7_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_5__5_  & (!\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9  # 
// !\u_fir|taps_5__7_ ))

	.dataa(\u_fir|taps_5__5_ ),
	.datab(\u_fir|taps_5__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z9 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N20
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52928 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_5__10_  $ \u_fir|taps_5__8_  $ !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z6 ) # GND
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5  = CARRY(\u_fir|taps_5__10_  & (\u_fir|taps_5__8_  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z6 ) # !\u_fir|taps_5__10_  & \u_fir|taps_5__8_  & 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z6 )

	.dataa(\u_fir|taps_5__10_ ),
	.datab(\u_fir|taps_5__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z6 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N4
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_5_filter_block_prod_mults28_0|d_5_  $ \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx39967z1  $ !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_5_  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx39967z1  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_5_  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx39967z1  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_5_ ),
	.datab(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx39967z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N8
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|tap_array_5_filter_block_prod_mults28_0|d_7_  $ !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|d_7_  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|tap_array_5_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N4
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52938 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_2_  = (\u_fir|taps_6__2_  $ \u_fir|taps_6__3_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z15 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14  = CARRY(\u_fir|taps_6__2_  & (\u_fir|taps_6__3_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z15 ) # !\u_fir|taps_6__2_  & \u_fir|taps_6__3_  & 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z15 )

	.dataa(\u_fir|taps_6__2_ ),
	.datab(\u_fir|taps_6__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z15 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_2_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52938 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N8
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52936 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_6__4_  $ \u_fir|taps_6__5_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z13 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12  = CARRY(\u_fir|taps_6__4_  & (\u_fir|taps_6__5_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z13 ) # !\u_fir|taps_6__4_  & \u_fir|taps_6__5_  & 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z13 )

	.dataa(\u_fir|taps_6__4_ ),
	.datab(\u_fir|taps_6__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z13 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52936 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N10
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52935 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_6__6_  & (\u_fir|taps_6__5_  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12  & VCC # !\u_fir|taps_6__5_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12 ) # 
// !\u_fir|taps_6__6_  & (\u_fir|taps_6__5_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12  # !\u_fir|taps_6__5_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12  # GND))
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z11  = CARRY(\u_fir|taps_6__6_  & !\u_fir|taps_6__5_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12  # !\u_fir|taps_6__6_  & (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12  
// # !\u_fir|taps_6__5_ ))

	.dataa(\u_fir|taps_6__6_ ),
	.datab(\u_fir|taps_6__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z12 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52935 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N12
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52934 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_6__6_  $ \u_fir|taps_6__7_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z11 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10  = CARRY(\u_fir|taps_6__6_  & (\u_fir|taps_6__7_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z11 ) # !\u_fir|taps_6__6_  & \u_fir|taps_6__7_  & 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z11 )

	.dataa(\u_fir|taps_6__6_ ),
	.datab(\u_fir|taps_6__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z11 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52934 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N18
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52931 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_6__9_  & (\u_fir|taps_6__10_  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8  & VCC # !\u_fir|taps_6__10_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8 ) # 
// !\u_fir|taps_6__9_  & (\u_fir|taps_6__10_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8  # !\u_fir|taps_6__10_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8  # GND))
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z7  = CARRY(\u_fir|taps_6__9_  & !\u_fir|taps_6__10_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8  # !\u_fir|taps_6__9_  & (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8  # 
// !\u_fir|taps_6__10_ ))

	.dataa(\u_fir|taps_6__9_ ),
	.datab(\u_fir|taps_6__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N6
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52947 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_3__dup_193  = \u_fir|tap_array_6_filter_block_prod_mults28_0|d_5_  & (\u_fir|taps_6__3_  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24  & VCC # !\u_fir|taps_6__3_  & 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24 ) # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_5_  & (\u_fir|taps_6__3_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24  # !\u_fir|taps_6__3_  & 
// (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24  # GND))
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z23  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_5_  & !\u_fir|taps_6__3_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24  # 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_5_  & (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24  # !\u_fir|taps_6__3_ ))

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_5_ ),
	.datab(\u_fir|taps_6__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_3__dup_193 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z23 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52947 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52947 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N8
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52946 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_4__dup_192  = (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6_  $ \u_fir|taps_6__4_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z23 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6_  & (\u_fir|taps_6__4_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z23 ) # 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6_  & \u_fir|taps_6__4_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z23 )

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6_ ),
	.datab(\u_fir|taps_6__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z23 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4__dup_192 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52946 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52946 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N12
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52944 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_6__dup_190  = (\u_fir|taps_6__6_  $ \u_fir|tap_array_6_filter_block_prod_mults28_0|d_8_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z21 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20  = CARRY(\u_fir|taps_6__6_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_8_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z21 ) # !\u_fir|taps_6__6_  & 
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z21 )

	.dataa(\u_fir|taps_6__6_ ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z21 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6__dup_190 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52944 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52944 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N16
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52942 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_8__dup_188  = (\u_fir|taps_6__8_  $ \u_fir|tap_array_6_filter_block_prod_mults28_0|d_10_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z19 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18  = CARRY(\u_fir|taps_6__8_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z19 ) # !\u_fir|taps_6__8_  & 
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z19 )

	.dataa(\u_fir|taps_6__8_ ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z19 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_8__dup_188 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52942 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52942 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N0
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_6_filter_block_prod_mults28_0|d_3__dup_193  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx37973z1  $ VCC) # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_3__dup_193 
//  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx37973z1  & VCC
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_3__dup_193  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx37973z1 )

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_3__dup_193 ),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx37973z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N2
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_6_filter_block_prod_mults28_0|d_4__dup_192  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4__dup_192  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1  & 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4__dup_192  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46  
// # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4__dup_192  & (!\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1 ))

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4__dup_192 ),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N6
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_6_filter_block_prod_mults28_0|d_6__dup_190  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6__dup_190  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1  & 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6__dup_190  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40  
// # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6__dup_190  & (!\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1 ))

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_6__dup_190 ),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N8
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|tap_array_6_filter_block_prod_mults28_0|d_7__dup_189  $ !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7__dup_189  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z37 ) 
// # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|tap_array_6_filter_block_prod_mults28_0|d_7__dup_189  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7__dup_189 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N10
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52931 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_7__6_  & (\u_fir|taps_7__5_  & \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9  & VCC # !\u_fir|taps_7__5_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9 ) # 
// !\u_fir|taps_7__6_  & (\u_fir|taps_7__5_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_7__5_  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9  # GND))
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z8  = CARRY(\u_fir|taps_7__6_  & !\u_fir|taps_7__5_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_7__6_  & (!\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9  # 
// !\u_fir|taps_7__5_ ))

	.dataa(\u_fir|taps_7__6_ ),
	.datab(\u_fir|taps_7__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N14
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52929 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_7__7_  & (\u_fir|taps_7__8_  & \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7  & VCC # !\u_fir|taps_7__8_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7 ) # 
// !\u_fir|taps_7__7_  & (\u_fir|taps_7__8_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_7__8_  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7  # GND))
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z6  = CARRY(\u_fir|taps_7__7_  & !\u_fir|taps_7__8_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_7__7_  & (!\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7  # 
// !\u_fir|taps_7__8_ ))

	.dataa(\u_fir|taps_7__7_ ),
	.datab(\u_fir|taps_7__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N16
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52928 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_7__9_  $ \u_fir|taps_7__8_  $ !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z6 ) # GND
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5  = CARRY(\u_fir|taps_7__9_  & (\u_fir|taps_7__8_  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z6 ) # !\u_fir|taps_7__9_  & \u_fir|taps_7__8_  & 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z6 )

	.dataa(\u_fir|taps_7__9_ ),
	.datab(\u_fir|taps_7__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z6 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N0
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_3_  $ VCC) # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx37973z1  & 
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_3_  & VCC
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|tap_array_7_filter_block_prod_mults28_0|d_3_ )

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N2
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_  & 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_ ))

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N4
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_5_  $ \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx39967z1  $ !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_5_  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx39967z1  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_5_  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx39967z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_5_ ),
	.datab(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx39967z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N8
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|tap_array_7_filter_block_prod_mults28_0|d_7_  $ !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_7_  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|tap_array_7_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N10
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_7_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_8_  & (!\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_8_ ),
	.datab(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N16
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52930 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_8__7_  $ \u_fir|taps_8__6_  $ !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z8 ) # GND
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7  = CARRY(\u_fir|taps_8__7_  & (\u_fir|taps_8__6_  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z8 ) # !\u_fir|taps_8__7_  & \u_fir|taps_8__6_  & 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z8 )

	.dataa(\u_fir|taps_8__7_ ),
	.datab(\u_fir|taps_8__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z8 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N2
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_  & 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_ ))

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N4
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|tap_array_8_filter_block_prod_mults28_0|d_5_  $ !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_5_  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|tap_array_8_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N8
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|tap_array_8_filter_block_prod_mults28_0|d_7_  $ !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_7_  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|tap_array_8_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52933 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_9__4_  & (\u_fir|taps_9__3_  & \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11  & VCC # !\u_fir|taps_9__3_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11 ) # 
// !\u_fir|taps_9__4_  & (\u_fir|taps_9__3_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_9__3_  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11  # GND))
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z10  = CARRY(\u_fir|taps_9__4_  & !\u_fir|taps_9__3_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_9__4_  & (!\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11  # 
// !\u_fir|taps_9__3_ ))

	.dataa(\u_fir|taps_9__4_ ),
	.datab(\u_fir|taps_9__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52930 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_9__7_  $ \u_fir|taps_9__6_  $ !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z8 ) # GND
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7  = CARRY(\u_fir|taps_9__7_  & (\u_fir|taps_9__6_  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z8 ) # !\u_fir|taps_9__7_  & \u_fir|taps_9__6_  & 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z8 )

	.dataa(\u_fir|taps_9__7_ ),
	.datab(\u_fir|taps_9__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z8 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52928 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_9__9_  $ \u_fir|taps_9__8_  $ !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z6 ) # GND
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5  = CARRY(\u_fir|taps_9__9_  & (\u_fir|taps_9__8_  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z6 ) # !\u_fir|taps_9__9_  & \u_fir|taps_9__8_  & 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z6 )

	.dataa(\u_fir|taps_9__9_ ),
	.datab(\u_fir|taps_9__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z6 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_  & 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_ ))

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|tap_array_9_filter_block_prod_mults28_0|d_5_  $ !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|d_5_  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|tap_array_9_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52933 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_10__4_  & (\u_fir|taps_10__3_  & \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11  & VCC # !\u_fir|taps_10__3_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11 ) # 
// !\u_fir|taps_10__4_  & (\u_fir|taps_10__3_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_10__3_  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11  # GND))
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z10  = CARRY(\u_fir|taps_10__4_  & !\u_fir|taps_10__3_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_10__4_  & 
// (!\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_10__3_ ))

	.dataa(\u_fir|taps_10__4_ ),
	.datab(\u_fir|taps_10__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52930 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_10__7_  $ \u_fir|taps_10__6_  $ !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z8 ) # GND
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7  = CARRY(\u_fir|taps_10__7_  & (\u_fir|taps_10__6_  # !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z8 ) # !\u_fir|taps_10__7_  & \u_fir|taps_10__6_  & 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z8 )

	.dataa(\u_fir|taps_10__7_ ),
	.datab(\u_fir|taps_10__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z8 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52929 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_10__7_  & (\u_fir|taps_10__8_  & \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7  & VCC # !\u_fir|taps_10__8_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7 ) # 
// !\u_fir|taps_10__7_  & (\u_fir|taps_10__8_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_10__8_  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7  # GND))
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z6  = CARRY(\u_fir|taps_10__7_  & !\u_fir|taps_10__8_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_10__7_  & (!\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7  
// # !\u_fir|taps_10__8_ ))

	.dataa(\u_fir|taps_10__7_ ),
	.datab(\u_fir|taps_10__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z7 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52928 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_10__9_  $ \u_fir|taps_10__8_  $ !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z6 ) # GND
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5  = CARRY(\u_fir|taps_10__9_  & (\u_fir|taps_10__8_  # !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z6 ) # !\u_fir|taps_10__9_  & \u_fir|taps_10__8_  & 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z6 )

	.dataa(\u_fir|taps_10__9_ ),
	.datab(\u_fir|taps_10__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z6 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_10_filter_block_prod_mults28_0|d_3_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx37973z1  $ VCC) # !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_3_  & 
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx37973z1  & VCC
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_3_  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx37973z1 )

	.dataa(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_3_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx37973z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_  & \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_  & 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_ ))

	.dataa(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|tap_array_10_filter_block_prod_mults28_0|d_5_  $ !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|d_5_  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|tap_array_10_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_10_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1  & \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1  & 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_6_  & (!\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1 ))

	.dataa(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_6_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_10_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_8_  & (!\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_8_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52929 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_11__8_  & (\u_fir|taps_11__7_  & \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7  & VCC # !\u_fir|taps_11__7_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7 ) # 
// !\u_fir|taps_11__8_  & (\u_fir|taps_11__7_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_11__7_  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7  # GND))
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z6  = CARRY(\u_fir|taps_11__8_  & !\u_fir|taps_11__7_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_11__8_  & (!\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7  
// # !\u_fir|taps_11__7_ ))

	.dataa(\u_fir|taps_11__8_ ),
	.datab(\u_fir|taps_11__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_3_  $ VCC) # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx37973z1  & 
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_3_  & VCC
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|tap_array_11_filter_block_prod_mults28_0|d_3_ )

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_  & 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_ ))

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_  & 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx40964z1  & (!\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_ ))

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx40964z1 ),
	.datab(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52938 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_2_  = (\u_fir|taps_12__2_  $ \u_fir|taps_12__3_  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z15 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14  = CARRY(\u_fir|taps_12__2_  & (\u_fir|taps_12__3_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z15 ) # !\u_fir|taps_12__2_  & \u_fir|taps_12__3_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z15 )

	.dataa(\u_fir|taps_12__2_ ),
	.datab(\u_fir|taps_12__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z15 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_2_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52938 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52937 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_12__4_  & (\u_fir|taps_12__3_  & \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14  & VCC # !\u_fir|taps_12__3_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14 ) # 
// !\u_fir|taps_12__4_  & (\u_fir|taps_12__3_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14  # !\u_fir|taps_12__3_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14  # GND))
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z13  = CARRY(\u_fir|taps_12__4_  & !\u_fir|taps_12__3_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14  # !\u_fir|taps_12__4_  & 
// (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14  # !\u_fir|taps_12__3_ ))

	.dataa(\u_fir|taps_12__4_ ),
	.datab(\u_fir|taps_12__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z14 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52937 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52933 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_12__7_  & (\u_fir|taps_12__8_  & \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10  & VCC # !\u_fir|taps_12__8_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10 ) # 
// !\u_fir|taps_12__7_  & (\u_fir|taps_12__8_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10  # !\u_fir|taps_12__8_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10  # GND))
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z9  = CARRY(\u_fir|taps_12__7_  & !\u_fir|taps_12__8_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10  # !\u_fir|taps_12__7_  & 
// (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10  # !\u_fir|taps_12__8_ ))

	.dataa(\u_fir|taps_12__7_ ),
	.datab(\u_fir|taps_12__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52932 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_12__9_  $ \u_fir|taps_12__8_  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z9 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8  = CARRY(\u_fir|taps_12__9_  & (\u_fir|taps_12__8_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z9 ) # !\u_fir|taps_12__9_  & \u_fir|taps_12__8_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z9 )

	.dataa(\u_fir|taps_12__9_ ),
	.datab(\u_fir|taps_12__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z9 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52930 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_12__15_  $ \u_fir|taps_12__10_  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z7 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z6  = CARRY(\u_fir|taps_12__15_  & (\u_fir|taps_12__10_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z7 ) # !\u_fir|taps_12__15_  & \u_fir|taps_12__10_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z7 )

	.dataa(\u_fir|taps_12__15_ ),
	.datab(\u_fir|taps_12__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z7 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52945 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_5__dup_191  = \u_fir|tap_array_12_filter_block_prod_mults28_0|d_7_  & (\u_fir|taps_12__5_  & \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22  & VCC # !\u_fir|taps_12__5_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22 ) # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7_  & (\u_fir|taps_12__5_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22  # !\u_fir|taps_12__5_  & 
// (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22  # GND))
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z21  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7_  & !\u_fir|taps_12__5_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22  # 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7_  & (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22  # !\u_fir|taps_12__5_ ))

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|taps_12__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5__dup_191 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z21 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52945 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52945 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52943 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_7__dup_189  = \u_fir|taps_12__7_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_  & \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20  & VCC # 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20 ) # !\u_fir|taps_12__7_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20  # GND))
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z19  = CARRY(\u_fir|taps_12__7_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20  # !\u_fir|taps_12__7_  & 
// (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_ ))

	.dataa(\u_fir|taps_12__7_ ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7__dup_189 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52943 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52943 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52942 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_8__dup_188  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10_  $ \u_fir|taps_12__8_  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z19 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10_  & (\u_fir|taps_12__8_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z19 ) # 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10_  & \u_fir|taps_12__8_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z19 )

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|taps_12__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z19 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8__dup_188 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52942 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52942 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5__dup_191  $ \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx39967z1  $ !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z43 ) # 
// GND
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5__dup_191  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx39967z1  # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z43 ) # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5__dup_191  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx39967z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5__dup_191 ),
	.datab(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx39967z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40  & 
// VCC # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx40964z1  & 
// (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40  
// # GND))
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190  & 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx40964z1  & (!\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190 
// ))

	.dataa(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx40964z1 ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52933 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_13__3_  & (\u_fir|taps_13__5_  & \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11  & VCC # !\u_fir|taps_13__5_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11 ) # 
// !\u_fir|taps_13__3_  & (\u_fir|taps_13__5_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_13__5_  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11  # GND))
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z10  = CARRY(\u_fir|taps_13__3_  & !\u_fir|taps_13__5_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_13__3_  & 
// (!\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_13__5_ ))

	.dataa(\u_fir|taps_13__3_ ),
	.datab(\u_fir|taps_13__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52932 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_13__6_  $ \u_fir|taps_13__4_  $ !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z10 ) # GND
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9  = CARRY(\u_fir|taps_13__6_  & (\u_fir|taps_13__4_  # !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z10 ) # !\u_fir|taps_13__6_  & \u_fir|taps_13__4_  & 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z10 )

	.dataa(\u_fir|taps_13__6_ ),
	.datab(\u_fir|taps_13__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z10 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52929 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_13__9_  & (\u_fir|taps_13__7_  & \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7  & VCC # !\u_fir|taps_13__7_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7 ) # 
// !\u_fir|taps_13__9_  & (\u_fir|taps_13__7_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_13__7_  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7  # GND))
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z6  = CARRY(\u_fir|taps_13__9_  & !\u_fir|taps_13__7_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_13__9_  & (!\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7  
// # !\u_fir|taps_13__7_ ))

	.dataa(\u_fir|taps_13__9_ ),
	.datab(\u_fir|taps_13__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52928 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_13__10_  $ \u_fir|taps_13__8_  $ !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z6 ) # GND
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5  = CARRY(\u_fir|taps_13__10_  & (\u_fir|taps_13__8_  # !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z6 ) # !\u_fir|taps_13__10_  & \u_fir|taps_13__8_  & 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z6 )

	.dataa(\u_fir|taps_13__10_ ),
	.datab(\u_fir|taps_13__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z6 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_13_filter_block_prod_mults28_0|d_3_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx37973z1  $ VCC) # !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_3_  & 
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx37973z1  & VCC
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_3_  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx37973z1 )

	.dataa(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_3_ ),
	.datab(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx37973z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_13_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1  & \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1  & 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_4_  & (!\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1 ))

	.dataa(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_4_ ),
	.datab(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|tap_array_13_filter_block_prod_mults28_0|d_5_  $ !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|d_5_  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|tap_array_13_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_13_filter_block_prod_mults28_0|d_7_  $ \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx41961z1  $ !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx41961z1  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_7_  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx41961z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx41961z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|taps_14__4_  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46  & VCC # !\u_fir|taps_14__4_  & 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|taps_14__4_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|taps_14__4_  & 
// (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|taps_14__4_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|taps_14__4_ ))

	.dataa(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|taps_14__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|taps_14__6_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|taps_14__6_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1  & 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|taps_14__6_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|taps_14__6_  & 
// (!\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1 ))

	.dataa(\u_fir|taps_14__6_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y12_N26
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52935 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_15__3_  & (\u_fir|taps_15__6_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13  # !\u_fir|taps_15__6_  & \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13  & VCC) # 
// !\u_fir|taps_15__3_  & (\u_fir|taps_15__6_  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13  # GND) # !\u_fir|taps_15__6_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13 )
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z12  = CARRY(\u_fir|taps_15__3_  & \u_fir|taps_15__6_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13  # !\u_fir|taps_15__3_  & (\u_fir|taps_15__6_  # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13 ))

	.dataa(\u_fir|taps_15__3_ ),
	.datab(\u_fir|taps_15__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52935 .lut_mask = 16'h694D;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y12_N30
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52933 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_15__5_  & (\u_fir|taps_15__8_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11  # !\u_fir|taps_15__8_  & \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11  & VCC) # 
// !\u_fir|taps_15__5_  & (\u_fir|taps_15__8_  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11  # GND) # !\u_fir|taps_15__8_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11 )
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z10  = CARRY(\u_fir|taps_15__5_  & \u_fir|taps_15__8_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11  # !\u_fir|taps_15__5_  & (\u_fir|taps_15__8_  # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11 ))

	.dataa(\u_fir|taps_15__5_ ),
	.datab(\u_fir|taps_15__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52933 .lut_mask = 16'h694D;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52931 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_15__10_  & (\u_fir|taps_15__7_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9  # !\u_fir|taps_15__7_  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9  # GND)) 
// # !\u_fir|taps_15__10_  & (\u_fir|taps_15__7_  & \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9  & VCC # !\u_fir|taps_15__7_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9 )
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z8  = CARRY(\u_fir|taps_15__10_  & (!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9  # !\u_fir|taps_15__7_ ) # !\u_fir|taps_15__10_  & !\u_fir|taps_15__7_  & 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9 )

	.dataa(\u_fir|taps_15__10_ ),
	.datab(\u_fir|taps_15__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52931 .lut_mask = 16'h692B;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52930 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_15__8_  $ \u_fir|taps_15__15_  $ \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z8 ) # GND
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7  = CARRY(\u_fir|taps_15__8_  & (!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z8  # !\u_fir|taps_15__15_ ) # !\u_fir|taps_15__8_  & !\u_fir|taps_15__15_  & 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z8 )

	.dataa(\u_fir|taps_15__8_ ),
	.datab(\u_fir|taps_15__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z8 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52930 .lut_mask = 16'h962B;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_15_filter_block_prod_mults28_0|d_5_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx37973z1  $ VCC) # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_5_  & 
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx37973z1  & VCC
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_5_  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx37973z1 )

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_5_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx37973z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_  & \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_  & 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_ ))

	.dataa(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_7_  $ \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx39967z1  $ !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx39967z1  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_7_  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx39967z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx39967z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_9_  $ \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx41961z1  $ !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_9_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx41961z1  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_9_  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx41961z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_9_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx41961z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_15_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_10_  & (!\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X44_Y14_N17
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__9_ ));

// atom is at LCCOMB_X44_Y14_N14
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52929 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_16__7_  & (\u_fir|taps_16__8_  & \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7  & VCC # !\u_fir|taps_16__8_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7 ) # 
// !\u_fir|taps_16__7_  & (\u_fir|taps_16__8_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7  # !\u_fir|taps_16__8_  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7  # GND))
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z6  = CARRY(\u_fir|taps_16__7_  & !\u_fir|taps_16__8_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7  # !\u_fir|taps_16__7_  & (!\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7  
// # !\u_fir|taps_16__8_ ))

	.dataa(\u_fir|taps_16__7_ ),
	.datab(\u_fir|taps_16__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N0
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|d_4_  $ VCC) # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx37973z1  & 
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_4_  & VCC
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|tap_array_16_filter_block_prod_mults28_0|d_4_ )

	.dataa(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N2
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_  & 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_ ))

	.dataa(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N4
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|tap_array_16_filter_block_prod_mults28_0|d_6_  $ !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|d_6_  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|tap_array_16_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N8
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|tap_array_16_filter_block_prod_mults28_0|d_8_  $ !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|d_8_  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|tap_array_16_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N10
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_  & 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx42958z1  & (!\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_ ))

	.dataa(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx42958z1 ),
	.datab(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X43_Y14_N17
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_7_ ));

// atom is at LCFF_X43_Y14_N21
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_9_ ));

// atom is at LCFF_X43_Y14_N13
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_5_ ));

// atom is at LCFF_X43_Y14_N9
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_3_ ));

// atom is at LCCOMB_X43_Y14_N14
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52932 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_6_  = (\u_fir|tap_array_17_filter_block_tap_next_9_  $ \u_fir|tap_array_17_filter_block_tap_next_6_  $ !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z10 ) # GND
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_9_  & (\u_fir|tap_array_17_filter_block_tap_next_6_  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z10 ) # 
// !\u_fir|tap_array_17_filter_block_tap_next_9_  & \u_fir|tap_array_17_filter_block_tap_next_6_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z10 )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_9_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z10 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N0
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_3_  $ VCC) # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx37973z1  & 
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_3_  & VCC
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|tap_array_17_filter_block_prod_mults28_0|d_3_ )

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N2
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_  & \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_  & 
// !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_ ))

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N8
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|tap_array_17_filter_block_prod_mults28_0|d_7_  $ !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_7_  # !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|tap_array_17_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N10
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_  & \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_  & 
// !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx42958z1  & (!\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_ ))

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx42958z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N18
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52929 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_1__9_  & (\u_fir|taps_1__15_  & \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7  & VCC # !\u_fir|taps_1__15_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7 ) # 
// !\u_fir|taps_1__9_  & (\u_fir|taps_1__15_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7  # !\u_fir|taps_1__15_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7  # GND))
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z6  = CARRY(\u_fir|taps_1__9_  & !\u_fir|taps_1__15_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7  # !\u_fir|taps_1__9_  & (!\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7  # 
// !\u_fir|taps_1__15_ ))

	.dataa(\u_fir|taps_1__9_ ),
	.datab(\u_fir|taps_1__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z7 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N20
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52926 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_2__15_  $ \u_fir|taps_2__10_  $ !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z4 ) # GND
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z3  = CARRY(\u_fir|taps_2__15_  & (\u_fir|taps_2__10_  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z4 ) # !\u_fir|taps_2__15_  & \u_fir|taps_2__10_  & 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z4 )

	.dataa(\u_fir|taps_2__15_ ),
	.datab(\u_fir|taps_2__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z4 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N12
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_2_filter_block_prod_mults28_0|d_10_  $ \u_fir|tap_array_1_filter_block_prod_mults28_0|d_9_  $ !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_9_  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_10_  & \u_fir|tap_array_1_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N6
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52929 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_11_  = \u_fir|taps_3__9_  & (\u_fir|taps_3__15_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7  # !\u_fir|taps_3__15_  & \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7  & VCC) # 
// !\u_fir|taps_3__9_  & (\u_fir|taps_3__15_  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7  # GND) # !\u_fir|taps_3__15_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7 )
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z6  = CARRY(\u_fir|taps_3__9_  & \u_fir|taps_3__15_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7  # !\u_fir|taps_3__9_  & (\u_fir|taps_3__15_  # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7 ))

	.dataa(\u_fir|taps_3__9_ ),
	.datab(\u_fir|taps_3__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z7 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52929 .lut_mask = 16'h694D;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N12
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_11_  $ \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx43955z1  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_11_ ),
	.datab(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N12
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|taps_4__9_  $ \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|taps_4__9_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx43955z1  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z31 ) # !\u_fir|taps_4__9_  & 
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|taps_4__9_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N22
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52927 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_5__15_  & (\u_fir|taps_5__9_  & \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5  & VCC # !\u_fir|taps_5__9_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5 ) # 
// !\u_fir|taps_5__15_  & (\u_fir|taps_5__9_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_5__9_  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5  # GND))
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z4  = CARRY(\u_fir|taps_5__15_  & !\u_fir|taps_5__9_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_5__15_  & (!\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5  # 
// !\u_fir|taps_5__9_ ))

	.dataa(\u_fir|taps_5__15_ ),
	.datab(\u_fir|taps_5__9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z5 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N12
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx43955z1  $ \u_fir|tap_array_5_filter_block_prod_mults28_0|d_9_  $ !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx43955z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|d_9_  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx43955z1  & \u_fir|tap_array_5_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx43955z1 ),
	.datab(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N22
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52929 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z6 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|b_10_  = CARRY(\u_fir|taps_6__15_ )

	.dataa(\u_fir|taps_6__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z6 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|b_10_ ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52929 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N18
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52941 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_9__dup_187  = \u_fir|taps_6__9_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18  & VCC # 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18 ) # !\u_fir|taps_6__9_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_  & 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18  # GND))
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z17  = CARRY(\u_fir|taps_6__9_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18  # !\u_fir|taps_6__9_  & 
// (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_ ))

	.dataa(\u_fir|taps_6__9_ ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z18 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9__dup_187 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z17 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52941 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52941 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N18
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52927 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_7__9_  & (\u_fir|taps_7__10_  & \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5  & VCC # !\u_fir|taps_7__10_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5 ) # 
// !\u_fir|taps_7__9_  & (\u_fir|taps_7__10_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_7__10_  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5  # GND))
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z4  = CARRY(\u_fir|taps_7__9_  & !\u_fir|taps_7__10_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_7__9_  & (!\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5  # 
// !\u_fir|taps_7__10_ ))

	.dataa(\u_fir|taps_7__9_ ),
	.datab(\u_fir|taps_7__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z5 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N22
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52927 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_8__9_  & (\u_fir|taps_8__10_  & \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5  & VCC # !\u_fir|taps_8__10_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5 ) # 
// !\u_fir|taps_8__9_  & (\u_fir|taps_8__10_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_8__10_  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5  # GND))
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z4  = CARRY(\u_fir|taps_8__9_  & !\u_fir|taps_8__10_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_8__9_  & (!\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5  # 
// !\u_fir|taps_8__10_ ))

	.dataa(\u_fir|taps_8__9_ ),
	.datab(\u_fir|taps_8__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N12
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_9_  $ \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_9_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx43955z1  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_9_  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_9_ ),
	.datab(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx43955z1  $ \u_fir|tap_array_9_filter_block_prod_mults28_0|d_9_  $ !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx43955z1  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|d_9_  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx43955z1  & \u_fir|tap_array_9_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx43955z1 ),
	.datab(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx43955z1  $ \u_fir|tap_array_10_filter_block_prod_mults28_0|d_9_  $ !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx43955z1  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|d_9_  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx43955z1  & \u_fir|tap_array_10_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx43955z1 ),
	.datab(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52941 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_9__dup_187  = \u_fir|taps_12__9_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18  & VCC # 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18 ) # !\u_fir|taps_12__9_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18  # GND))
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z17  = CARRY(\u_fir|taps_12__9_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18  # !\u_fir|taps_12__9_  & 
// (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_ ))

	.dataa(\u_fir|taps_12__9_ ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z18 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9__dup_187 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z17 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52941 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52941 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9__dup_187  $ \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z31 ) # 
// GND
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9__dup_187  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx43955z1  # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z31 ) # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9__dup_187  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9__dup_187 ),
	.datab(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52929 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_11_  = \u_fir|taps_15__15_  & (\u_fir|taps_15__9_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7  # !\u_fir|taps_15__9_  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7  # GND)) 
// # !\u_fir|taps_15__15_  & (\u_fir|taps_15__9_  & \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7  & VCC # !\u_fir|taps_15__9_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7 )
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z6  = CARRY(\u_fir|taps_15__15_  & (!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7  # !\u_fir|taps_15__9_ ) # !\u_fir|taps_15__15_  & !\u_fir|taps_15__9_  & 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7 )

	.dataa(\u_fir|taps_15__15_ ),
	.datab(\u_fir|taps_15__9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z7 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52929 .lut_mask = 16'h692B;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N20
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52926 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_16__15_  $ \u_fir|taps_16__10_  $ !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z4 ) # GND
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z3  = CARRY(\u_fir|taps_16__15_  & (\u_fir|taps_16__10_  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z4 ) # !\u_fir|taps_16__15_  & \u_fir|taps_16__10_  & 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z4 )

	.dataa(\u_fir|taps_16__15_ ),
	.datab(\u_fir|taps_16__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z4 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N12
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_16_filter_block_prod_mults28_0|d_10_  $ \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx43955z1  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_10_  & \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N20
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52928 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_1__10_  $ \u_fir|taps_1__15_  $ !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z6 ) # GND
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z5  = CARRY(\u_fir|taps_1__10_  & (\u_fir|taps_1__15_  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z6 ) # !\u_fir|taps_1__10_  & \u_fir|taps_1__15_  & 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z6 )

	.dataa(\u_fir|taps_1__10_ ),
	.datab(\u_fir|taps_1__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z6 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N22
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52925 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z3 ) # GND
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z2  = CARRY(\u_fir|taps_2__15_ )

	.dataa(\u_fir|taps_2__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z3 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N14
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_1_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_  & 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_10_  & (!\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_ ))

	.dataa(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N8
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52928 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_  = (\u_fir|taps_3__10_  $ \u_fir|taps_3__15_  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z6 ) # GND
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z5  = CARRY(\u_fir|taps_3__10_  & (!\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z6  # !\u_fir|taps_3__15_ ) # !\u_fir|taps_3__10_  & !\u_fir|taps_3__15_  & 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z6 )

	.dataa(\u_fir|taps_3__10_ ),
	.datab(\u_fir|taps_3__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z6 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52928 .lut_mask = 16'h962B;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N14
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_  & \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_  & 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx44952z1  & (!\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_ ))

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx44952z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_12_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N14
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|taps_4__10_  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28  & VCC # !\u_fir|taps_4__10_  & 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|taps_4__10_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|taps_4__10_  & 
// (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|taps_4__10_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx44952z1  & (!\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|taps_4__10_ ))

	.dataa(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx44952z1 ),
	.datab(\u_fir|taps_4__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N24
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52926 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_5__10_  $ \u_fir|taps_5__15_  $ !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z4 ) # GND
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z3  = CARRY(\u_fir|taps_5__10_  & (\u_fir|taps_5__15_  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z4 ) # !\u_fir|taps_5__10_  & \u_fir|taps_5__15_  & 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z4 )

	.dataa(\u_fir|taps_5__10_ ),
	.datab(\u_fir|taps_5__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z4 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N14
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_  & 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx44952z1  & (!\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_ ))

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx44952z1 ),
	.datab(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N24
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|ix10225z52928 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z5  = \u_fir|tap_array_6_filter_block_prod_mults28_0|b_10_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|b_10_ ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z5 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|ix10225z52928 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|ix10225z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N20
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52926 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_7__15_  $ \u_fir|taps_7__10_  $ !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z4 ) # GND
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z3  = CARRY(\u_fir|taps_7__15_  & (\u_fir|taps_7__10_  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z4 ) # !\u_fir|taps_7__15_  & \u_fir|taps_7__10_  & 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z4 )

	.dataa(\u_fir|taps_7__15_ ),
	.datab(\u_fir|taps_7__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z4 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N14
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_7_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1  & 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_10_  & (!\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1 ))

	.dataa(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N24
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52926 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_8__15_  $ \u_fir|taps_8__10_  $ !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z4 ) # GND
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z3  = CARRY(\u_fir|taps_8__15_  & (\u_fir|taps_8__10_  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z4 ) # !\u_fir|taps_8__15_  & \u_fir|taps_8__10_  & 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z4 )

	.dataa(\u_fir|taps_8__15_ ),
	.datab(\u_fir|taps_8__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z4 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52926 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_9__15_  $ \u_fir|taps_9__10_  $ !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z4 ) # GND
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z3  = CARRY(\u_fir|taps_9__15_  & (\u_fir|taps_9__10_  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z4 ) # !\u_fir|taps_9__15_  & \u_fir|taps_9__10_  & 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z4 )

	.dataa(\u_fir|taps_9__15_ ),
	.datab(\u_fir|taps_9__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z4 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52926 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_10__15_  $ \u_fir|taps_10__10_  $ !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z4 ) # GND
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z3  = CARRY(\u_fir|taps_10__15_  & (\u_fir|taps_10__10_  # !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z4 ) # !\u_fir|taps_10__15_  & \u_fir|taps_10__10_  & 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z4 )

	.dataa(\u_fir|taps_10__15_ ),
	.datab(\u_fir|taps_10__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z4 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_10_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1  & \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1  & 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_10_  & (!\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1 ))

	.dataa(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52927 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_10__dup_186  = (\u_fir|taps_12__10_  $ \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z5  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z17 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z4  = CARRY(\u_fir|taps_12__10_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z5  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z17 ) # !\u_fir|taps_12__10_  & 
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z5  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z17 )

	.dataa(\u_fir|taps_12__10_ ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z5 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z17 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10__dup_186 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52926 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_13__10_  $ \u_fir|taps_13__15_  $ !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z4 ) # GND
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z3  = CARRY(\u_fir|taps_13__10_  & (\u_fir|taps_13__15_  # !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z4 ) # !\u_fir|taps_13__10_  & \u_fir|taps_13__15_  & 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z4 )

	.dataa(\u_fir|taps_13__10_ ),
	.datab(\u_fir|taps_13__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z4 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_13_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1  & \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1  & 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_10_  & (!\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1 ))

	.dataa(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52928 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_12_  = (\u_fir|taps_15__10_  $ \u_fir|taps_15__15_  $ \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z6 ) # GND
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z5  = CARRY(\u_fir|taps_15__10_  & (!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z6  # !\u_fir|taps_15__15_ ) # !\u_fir|taps_15__10_  & !\u_fir|taps_15__15_  & 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z6 )

	.dataa(\u_fir|taps_15__10_ ),
	.datab(\u_fir|taps_15__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z6 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_12_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52928 .lut_mask = 16'h962B;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N22
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52925 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z3 ) # GND
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z2  = CARRY(\u_fir|taps_16__15_ )

	.dataa(\u_fir|taps_16__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z3 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N22
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52928 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_10_  = (\u_fir|tap_array_17_filter_block_tap_next_15_  $ \u_fir|tap_array_17_filter_block_tap_next_10_  $ !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z6 ) # GND
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z5  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_15_  & (\u_fir|tap_array_17_filter_block_tap_next_10_  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z6 ) # 
// !\u_fir|tap_array_17_filter_block_tap_next_15_  & \u_fir|tap_array_17_filter_block_tap_next_10_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z6 )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z6 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at M4K_X26_Y14
cycloneii_ram_block \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 (
	.portawe(gnd),
	.portaaddrstall(gnd),
	.portbrewe(vcc),
	.portbaddrstall(gnd),
	.clk0(\aud_adclrck_dup0~clkctrl_outclk ),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(12'b000000000000),
	.portaaddr({\u_sine_address_add9_0i1|nx45949z1 ,\u_sine_address_add9_0i1|nx44952z1 ,\u_sine_address_add9_0i1|nx43955z1 ,\u_sine_address_add9_0i1|nx42958z1 ,\u_sine_address_add9_0i1|nx41961z1 ,\u_sine_address_add9_0i1|nx40964z1 }),
	.portabyteenamasks(1'b1),
	.portbdatain(12'b000000000000),
	.portbaddr(6'b000000),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0_PORTADATAOUT_bus ),
	.portbdataout());
// synopsys translate_off
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .init_file = "u_sine_modgen_rom_ix21__altsyncram_12_6_64_2_0.hex";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .init_file_layout = "port_a";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .logical_ram_name = "altsyncram:u_sine_modgen_rom_ix21__ix62120z58996|altsyncram_0bk2:auto_generated|ALTSYNCRAM";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .operation_mode = "rom";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_address_width = 6;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_byte_enable_clear = "none";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_byte_enable_clock = "none";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_data_in_clear = "none";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_data_width = 12;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_last_address = 63;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 64;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_logical_ram_width = 12;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_write_enable_clear = "none";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_a_write_enable_clock = "none";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_b_address_width = 6;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .port_b_data_width = 12;
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .ram_block_type = "M4K";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .safe_write = "err_on_2clk";
defparam \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|ram_block1a0 .mem_init0 = 768'hF37E70DADCF0C3AB8EAECA579D09598F189B85882780980080982785889B8F19599D0A57AECB11C3ACF0DADE70F370000C818F25230F3C54715135A862F6A670E7647A77D87F67FF7F67D87A776470E6A662F5A85134713C530F25218F0C8000;
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N22
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52927 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z5 ) # GND
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z4  = CARRY(\u_fir|taps_1__15_ )

	.dataa(vcc),
	.datab(\u_fir|taps_1__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z5 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52927 .lut_mask = 16'hF0CC;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N24
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52926 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_12_  = (\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z4 ) # GND
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z3  = CARRY(\u_fir|taps_1__15_ )

	.dataa(vcc),
	.datab(\u_fir|taps_1__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z4 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_12_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52926 .lut_mask = 16'hF0CC;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N24
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|ix8231z52923 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z1  = \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z2 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|ix8231z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|ix8231z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N16
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_11_  $ \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z1  $ !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z1  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z1  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_11_ ),
	.datab(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N18
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_1_filter_block_prod_mults28_0|d_12_  & (\u_fir|taps_2__15_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22  & VCC # !\u_fir|taps_2__15_  & 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_12_  & (\u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|taps_2__15_  & 
// (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_12_  & !\u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_12_  & (!\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|taps_2__15_ ))

	.dataa(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_12_ ),
	.datab(\u_fir|taps_2__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N10
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52927 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_13_  = !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z5 
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z4  = CARRY(!\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z5 )

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z5 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_13_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52927 .lut_mask = 16'h0F0F;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N12
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52926 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_  = \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z4  $ GND
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z3  = CARRY(!\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z4 )

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z4 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52926 .lut_mask = 16'hF00F;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N16
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|d_13_  $ !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_13_  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_3_filter_block_prod_mults28_0|d_13_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_13_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N18
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_  & \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_  & 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx46946z1  & (!\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_ ))

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx46946z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_14_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N16
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|taps_4__15_  $ \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx45949z1  $ !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|taps_4__15_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx45949z1  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z25 ) # !\u_fir|taps_4__15_  & 
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx45949z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|taps_4__15_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx45949z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N18
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|taps_4__15_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|taps_4__15_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|taps_4__15_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|taps_4__15_  & 
// (!\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|taps_4__15_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N26
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52925 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z3 ) # GND
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z2  = CARRY(\u_fir|taps_5__15_ )

	.dataa(\u_fir|taps_5__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z3 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N28
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|ix9228z52923 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1  = \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z2 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|ix9228z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|ix9228z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N16
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_5_filter_block_prod_mults28_0|d_11_  $ !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|d_11_  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_5_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N18
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1  & 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx46946z1  & (!\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1 ))

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx46946z1 ),
	.datab(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N22
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52926 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_11__dup_185  = (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z4 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z3  = CARRY(\u_fir|taps_6__15_ )

	.dataa(\u_fir|taps_6__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z4 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11__dup_185 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52926 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N24
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52925 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_  = (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z3 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z2  = CARRY(\u_fir|taps_6__15_ )

	.dataa(\u_fir|taps_6__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z3 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N16
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_6_filter_block_prod_mults28_0|d_11__dup_185  $ !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z25 ) # 
// GND
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11__dup_185  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z25 
// ) # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_6_filter_block_prod_mults28_0|d_11__dup_185  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_11__dup_185 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N18
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_  & 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx46946z1  & (!\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_ ))

	.dataa(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx46946z1 ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_12_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N22
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52925 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z3 ) # GND
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z2  = CARRY(\u_fir|taps_7__15_ )

	.dataa(\u_fir|taps_7__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z3 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N24
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|ix9228z52923 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z1  = \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z2 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|ix9228z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|ix9228z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N16
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_11_  $ \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx45949z1  $ !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx45949z1  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx45949z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_11_ ),
	.datab(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx45949z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N18
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z1  & (!\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z1 ),
	.datab(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N26
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52925 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z3 ) # GND
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z2  = CARRY(\u_fir|taps_8__15_ )

	.dataa(\u_fir|taps_8__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z3 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N28
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|ix9228z52923 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1  = \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z2 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|ix9228z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|ix9228z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N16
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_11_  $ \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx45949z1  $ !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx45949z1  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx45949z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_11_ ),
	.datab(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx45949z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N18
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1  & 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx46946z1  & (!\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1 ))

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx46946z1 ),
	.datab(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52925 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z3 ) # GND
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z2  = CARRY(\u_fir|taps_9__15_ )

	.dataa(\u_fir|taps_9__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z3 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_9_filter_block_prod_mults28_0|d_11_  $ \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx45949z1  $ !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx45949z1  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx45949z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_11_ ),
	.datab(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx45949z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1  & 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx46946z1  & (!\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1 ))

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx46946z1 ),
	.datab(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52925 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z3 ) # GND
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z2  = CARRY(\u_fir|taps_10__15_ )

	.dataa(\u_fir|taps_10__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z3 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|ix9228z52923 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z1  = \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z2 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|ix9228z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|ix9228z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_10_filter_block_prod_mults28_0|d_11_  $ !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|d_11_  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_10_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z1  & (!\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z1 ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52925 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z3 ) # GND
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z2  = CARRY(\u_fir|taps_11__15_ )

	.dataa(vcc),
	.datab(\u_fir|taps_11__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z3 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52925 .lut_mask = 16'hF0CC;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|ix9228z52923 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z1  = \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z2 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|ix9228z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|ix9228z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22  
// # !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z1  & (!\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z1 ),
	.datab(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52926 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_11__dup_185  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z4 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z3  = CARRY(\u_fir|taps_12__15_ )

	.dataa(vcc),
	.datab(\u_fir|taps_12__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z4 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11__dup_185 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52926 .lut_mask = 16'hF0CC;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52925 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z3 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z2  = CARRY(\u_fir|taps_12__15_ )

	.dataa(vcc),
	.datab(\u_fir|taps_12__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z3 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52925 .lut_mask = 16'hF0CC;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11__dup_185  $ \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx45949z1  $ !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z25 ) 
// # GND
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11__dup_185  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx45949z1  # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z25 ) # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11__dup_185  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx45949z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z25 
// )

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11__dup_185 ),
	.datab(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx45949z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52925 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z3 ) # GND
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z2  = CARRY(\u_fir|taps_13__15_ )

	.dataa(\u_fir|taps_13__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z3 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|ix9228z52923 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z1  = \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z2 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|ix9228z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|ix9228z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|taps_14__15_  $ \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx45949z1  $ !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx45949z1  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z25 ) # !\u_fir|taps_14__15_  & 
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx45949z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|taps_14__15_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx45949z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52926 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_14_  = \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z4  $ GND
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z3  = CARRY(!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z4 )

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z4 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_14_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52926 .lut_mask = 16'hF00F;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_15_filter_block_prod_mults28_0|d_13_  $ !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_13_  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_15_filter_block_prod_mults28_0|d_13_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_13_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N16
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z1  $ !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z1  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z25 ) 
// # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N26
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52926 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_12_  = (\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z4 ) # GND
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z3  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_15_ )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z4 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_12_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52926 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N26
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52925 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_  = (\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z3 ) # GND
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z2  = CARRY(\u_fir|taps_1__15_ )

	.dataa(vcc),
	.datab(\u_fir|taps_1__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z3 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52925 .lut_mask = 16'hF0CC;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N20
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_  $ \u_fir|taps_2__15_  $ !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_  & (\u_fir|taps_2__15_  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_  & \u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_ ),
	.datab(\u_fir|taps_2__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N14
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52925 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_  = !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z3 
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z2  = CARRY(!\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z3 )

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z3 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52925 .lut_mask = 16'h0F0F;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N20
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_  $ \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx62798z1  $ !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx62798z1  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx62798z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_ ),
	.datab(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx62798z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N20
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|taps_4__15_  $ \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx62798z1  $ !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|taps_4__15_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx62798z1  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z19 ) # !\u_fir|taps_4__15_  & 
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx62798z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|taps_4__15_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx62798z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N20
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx62798z1  $ \u_fir|taps_5__15_  $ !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx62798z1  & (\u_fir|taps_5__15_  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx62798z1  & \u_fir|taps_5__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx62798z1 ),
	.datab(\u_fir|taps_5__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N26
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|ix10225z52923 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z1  = \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z2 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|ix10225z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|ix10225z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N20
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx62798z1  $ \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z1  $ !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx62798z1  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z1  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx62798z1  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx62798z1 ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N20
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx62798z1  $ \u_fir|taps_7__15_  $ !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx62798z1  & (\u_fir|taps_7__15_  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx62798z1  & \u_fir|taps_7__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx62798z1 ),
	.datab(\u_fir|taps_7__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N20
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx62798z1  $ \u_fir|taps_8__15_  $ !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx62798z1  & (\u_fir|taps_8__15_  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx62798z1  & \u_fir|taps_8__15_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx62798z1 ),
	.datab(\u_fir|taps_8__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx62798z1  $ \u_fir|taps_9__15_  $ !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx62798z1  & (\u_fir|taps_9__15_  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx62798z1  & \u_fir|taps_9__15_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx62798z1 ),
	.datab(\u_fir|taps_9__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|taps_10__15_  $ \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx62798z1  $ !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|taps_10__15_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx62798z1  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z19 ) # !\u_fir|taps_10__15_  & 
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx62798z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|taps_10__15_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx62798z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx62798z1  $ \u_fir|taps_11__15_  $ !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx62798z1  & (\u_fir|taps_11__15_  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx62798z1  & \u_fir|taps_11__15_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx62798z1 ),
	.datab(\u_fir|taps_11__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N30
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|ix10225z52923 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z1  = \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z2 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|ix10225z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|ix10225z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z1  $ \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx62798z1  $ !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z19 ) # 
// GND
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z1  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx62798z1  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z19 
// ) # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z1  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx62798z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z1 ),
	.datab(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx62798z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52925 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_  = !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z3 
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z2  = CARRY(!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z3 )

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z3 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52925 .lut_mask = 16'h0F0F;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N20
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|taps_16__15_  $ \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx62798z1  $ !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx62798z1  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z19 ) # !\u_fir|taps_16__15_  & 
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx62798z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|taps_16__15_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx62798z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N28
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52925 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  = (\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z3 ) # GND
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z2  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_15_ )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z3 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z2 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52925 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N22
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_  & (\u_fir|taps_2__15_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16  & VCC # !\u_fir|taps_2__15_  & 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_  & (\u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_2__15_  & 
// (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_  & !\u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_  & (!\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_2__15_ ))

	.dataa(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_13_ ),
	.datab(\u_fir|taps_2__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N22
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1  & \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1  & 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_  & (!\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1 ))

	.dataa(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_15_ ),
	.datab(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx63795z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N22
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|taps_4__15_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|taps_4__15_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1  & 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|taps_4__15_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_4__15_  & 
// (!\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1 ))

	.dataa(\u_fir|taps_4__15_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx63795z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N22
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_5__15_  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16  & VCC # !\u_fir|taps_5__15_  & 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_5__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_5__15_  & 
// (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|taps_5__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx63795z1  & (!\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_5__15_ ))

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx63795z1 ),
	.datab(\u_fir|taps_5__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N22
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|taps_6__15_  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|taps_6__15_  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1  & 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|taps_6__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_6__15_  & 
// (!\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1 ))

	.dataa(\u_fir|taps_6__15_ ),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx63795z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N22
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_7__15_  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16  & VCC # !\u_fir|taps_7__15_  & 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_7__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_7__15_  & 
// (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|taps_7__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx63795z1  & (!\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_7__15_ ))

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx63795z1 ),
	.datab(\u_fir|taps_7__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N22
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|taps_8__15_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|taps_8__15_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1  & 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|taps_8__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_8__15_  & 
// (!\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1 ))

	.dataa(\u_fir|taps_8__15_ ),
	.datab(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx63795z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_9__15_  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16  & VCC # !\u_fir|taps_9__15_  & 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_9__15_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_9__15_  & 
// (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|taps_9__15_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx63795z1  & (!\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_9__15_ ))

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx63795z1 ),
	.datab(\u_fir|taps_9__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|taps_10__15_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1  & \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|taps_10__15_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1  & 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|taps_10__15_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_10__15_  & 
// (!\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1 ))

	.dataa(\u_fir|taps_10__15_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx63795z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_11__15_  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16  & VCC # !\u_fir|taps_11__15_  & 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_11__15_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_11__15_  & 
// (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|taps_11__15_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx63795z1  & (!\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_11__15_ ))

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx63795z1 ),
	.datab(\u_fir|taps_11__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_12__15_  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16  & VCC # !\u_fir|taps_12__15_  & 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_12__15_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_12__15_  & 
// (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|taps_12__15_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx63795z1  & (!\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_12__15_ ))

	.dataa(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx63795z1 ),
	.datab(\u_fir|taps_12__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_13__15_  & \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16  & VCC # !\u_fir|taps_13__15_  & 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|taps_13__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_13__15_  & 
// (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|taps_13__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx63795z1  & (!\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_13__15_ ))

	.dataa(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx63795z1 ),
	.datab(\u_fir|taps_13__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1  & 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|taps_14__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_14__15_  & 
// (!\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1 ))

	.dataa(\u_fir|taps_14__15_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx63795z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N22
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1  & 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|taps_16__15_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|taps_16__15_  & 
// (!\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1 ))

	.dataa(\u_fir|taps_16__15_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N28
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52923 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z1  = \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z2 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N24
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z1  $ \u_fir|taps_2__15_  $ !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z1  & (\u_fir|taps_2__15_  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z1  & \u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z1 ),
	.datab(\u_fir|taps_2__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N26
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx253z1  = \u_fir|taps_1__15_  & (\u_fir|taps_2__15_  & \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10 
// ) # !\u_fir|taps_1__15_  & (\u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_2__15_  & (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|taps_1__15_  & !\u_fir|taps_2__15_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_1__15_  & 
// (!\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_2__15_ ))

	.dataa(\u_fir|taps_1__15_ ),
	.datab(\u_fir|taps_2__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N16
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52923 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  = \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z2 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N24
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  $ !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N26
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  & \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10  & VCC # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  & 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1 ))

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N24
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|taps_4__15_  $ \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx64792z1  $ !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|taps_4__15_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx64792z1  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z13 ) # !\u_fir|taps_4__15_  & 
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx64792z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|taps_4__15_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx64792z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N26
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_4__15_  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_4__15_  & 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_4__15_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_4__15_  & 
// (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|taps_4__15_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_4__15_ ))

	.dataa(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|taps_4__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N24
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|taps_5__15_  $ !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|taps_5__15_  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|taps_5__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|taps_5__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N26
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_5__15_  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_5__15_  & 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_5__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_5__15_  & 
// (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|taps_5__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_5__15_ ))

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|taps_5__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N24
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|taps_6__15_  $ \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx64792z1  $ !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|taps_6__15_  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx64792z1  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z13 ) # !\u_fir|taps_6__15_  & 
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx64792z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|taps_6__15_ ),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx64792z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N26
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx253z1  = \u_fir|taps_6__15_  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10  & VCC # 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|taps_6__15_  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1  & 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|taps_6__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_6__15_  & 
// (!\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1 ))

	.dataa(\u_fir|taps_6__15_ ),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx253z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N24
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|taps_7__15_  $ !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|taps_7__15_  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|taps_7__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|taps_7__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N26
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_7__15_  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_7__15_  & 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_7__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_7__15_  & 
// (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|taps_7__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_7__15_ ))

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|taps_7__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N24
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|taps_8__15_  $ !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|taps_8__15_  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|taps_8__15_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|taps_8__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N26
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx253z1  = \u_fir|taps_8__15_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10  & VCC # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|taps_8__15_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1  & 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|taps_8__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_8__15_  & 
// (!\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1 ))

	.dataa(\u_fir|taps_8__15_ ),
	.datab(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx253z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|taps_9__15_  $ !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|taps_9__15_  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|taps_9__15_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|taps_9__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_9__15_  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_9__15_  & 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_9__15_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_9__15_  & 
// (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|taps_9__15_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_9__15_ ))

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|taps_9__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|taps_10__15_  $ \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx64792z1  $ !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|taps_10__15_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx64792z1  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z13 ) # !\u_fir|taps_10__15_  & 
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx64792z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|taps_10__15_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx64792z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_10__15_  & \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_10__15_  & 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_10__15_  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_10__15_  & 
// (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|taps_10__15_  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_10__15_ ))

	.dataa(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|taps_10__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|taps_11__15_  $ !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|taps_11__15_  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|taps_11__15_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|taps_11__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_11__15_  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_11__15_  & 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_11__15_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_11__15_  & 
// (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|taps_11__15_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_11__15_ ))

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|taps_11__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|taps_12__15_  $ !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|taps_12__15_  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|taps_12__15_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|taps_12__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_12__15_  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_12__15_  & 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_12__15_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_12__15_  & 
// (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|taps_12__15_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_12__15_ ))

	.dataa(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|taps_12__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|taps_13__15_  $ !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|taps_13__15_  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z13 ) # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|taps_13__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|taps_13__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_13__15_  & \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10  & VCC # !\u_fir|taps_13__15_  & 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|taps_13__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_13__15_  & 
// (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|taps_13__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_13__15_ ))

	.dataa(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|taps_13__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|taps_14__15_  $ \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx64792z1  $ !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx64792z1  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z13 ) # !\u_fir|taps_14__15_  & 
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx64792z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|taps_14__15_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx64792z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx253z1  = \u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10  & VCC # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1  & 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|taps_14__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_14__15_  & 
// (!\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1 ))

	.dataa(\u_fir|taps_14__15_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx253z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N30
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52923 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z1  = \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z2 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N28
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|taps_1__15_  $ \u_fir|taps_2__15_  $ !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|taps_1__15_  & (\u_fir|taps_2__15_  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z7 ) # !\u_fir|taps_1__15_  & \u_fir|taps_2__15_  & 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|taps_1__15_ ),
	.datab(\u_fir|taps_2__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N28
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx1250z1  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  $ !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx1250z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx1250z1  & \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx1250z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N28
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|taps_4__15_  $ \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx1250z1  $ !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|taps_4__15_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx1250z1  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z7 ) # !\u_fir|taps_4__15_  & 
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx1250z1  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|taps_4__15_ ),
	.datab(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx1250z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N28
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx1250z1  $ \u_fir|taps_5__15_  $ !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx1250z1  & (\u_fir|taps_5__15_  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx1250z1  & \u_fir|taps_5__15_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx1250z1 ),
	.datab(\u_fir|taps_5__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N28
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx1250z1  $ \u_fir|taps_6__15_  $ !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx1250z1  & (\u_fir|taps_6__15_  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx1250z1  & \u_fir|taps_6__15_  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx1250z1 ),
	.datab(\u_fir|taps_6__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N28
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx1250z1  $ \u_fir|taps_7__15_  $ !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx1250z1  & (\u_fir|taps_7__15_  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx1250z1  & \u_fir|taps_7__15_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx1250z1 ),
	.datab(\u_fir|taps_7__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N28
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx1250z1  $ \u_fir|taps_8__15_  $ !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx1250z1  & (\u_fir|taps_8__15_  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx1250z1  & \u_fir|taps_8__15_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx1250z1 ),
	.datab(\u_fir|taps_8__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|taps_9__15_  $ \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx1250z1  $ !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|taps_9__15_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx1250z1  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z7 ) # !\u_fir|taps_9__15_  & 
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx1250z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|taps_9__15_ ),
	.datab(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx1250z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|taps_10__15_  $ \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx1250z1  $ !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|taps_10__15_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx1250z1  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z7 ) # !\u_fir|taps_10__15_  & 
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx1250z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|taps_10__15_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx1250z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|taps_11__15_  $ \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx1250z1  $ !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|taps_11__15_  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx1250z1  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z7 ) # !\u_fir|taps_11__15_  & 
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx1250z1  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|taps_11__15_ ),
	.datab(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx1250z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx1250z1  $ \u_fir|taps_12__15_  $ !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx1250z1  & (\u_fir|taps_12__15_  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx1250z1  & \u_fir|taps_12__15_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx1250z1 ),
	.datab(\u_fir|taps_12__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx1250z1  $ \u_fir|taps_13__15_  $ !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx1250z1  & (\u_fir|taps_13__15_  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx1250z1  & \u_fir|taps_13__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx1250z1 ),
	.datab(\u_fir|taps_13__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|taps_14__15_  $ \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx1250z1  $ !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx1250z1  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z7 ) # !\u_fir|taps_14__15_  & 
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx1250z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|taps_14__15_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx1250z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx1250z1  $ \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  $ !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx1250z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx1250z1  & \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx1250z1 ),
	.datab(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N28
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|taps_16__15_  $ \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx1250z1  $ !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx1250z1  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z7 ) # !\u_fir|taps_16__15_  & 
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx1250z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|taps_16__15_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx1250z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N28
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52925 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx1250z1  = (\u_fir|tap_array_17_filter_block_tap_next_15_  $ \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx1250z1  $ !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z7 ) # GND
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z4  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_15_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx1250z1  # !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z7 ) # 
// !\u_fir|tap_array_17_filter_block_tap_next_15_  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx1250z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z7 )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datab(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx1250z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z7 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx1250z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52925 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N30
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|taps_1__15_  $ \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|taps_2__15_ 

	.dataa(\u_fir|taps_1__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_2__15_ ),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hA55A;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N30
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z1  $ \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1 

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z1 ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z1 ),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hA55A;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N30
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|taps_4__15_  $ \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(\u_fir|taps_4__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hA55A;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N30
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z1  $ \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|taps_5__15_ 

	.dataa(vcc),
	.datab(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z1 ),
	.datac(vcc),
	.datad(\u_fir|taps_5__15_ ),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hC33C;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N30
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z1  $ \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|taps_6__15_ 

	.dataa(vcc),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z1 ),
	.datac(vcc),
	.datad(\u_fir|taps_6__15_ ),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hC33C;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N30
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z1  $ \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|taps_7__15_ 

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z1 ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_7__15_ ),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hA55A;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N30
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z1  $ \u_fir|taps_8__15_  $ \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z4 

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z1 ),
	.datab(\u_fir|taps_8__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'h9696;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N30
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z1  $ \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|taps_9__15_ 

	.dataa(vcc),
	.datab(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z1 ),
	.datac(vcc),
	.datad(\u_fir|taps_9__15_ ),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hC33C;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N30
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|taps_10__15_  $ \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(\u_fir|taps_10__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hA55A;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N30
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|taps_11__15_  $ \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(vcc),
	.datab(\u_fir|taps_11__15_ ),
	.datac(vcc),
	.datad(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hC33C;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N30
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|taps_12__15_  $ \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(vcc),
	.datab(\u_fir|taps_12__15_ ),
	.datac(vcc),
	.datad(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hC33C;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N30
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|taps_13__15_  $ \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(vcc),
	.datab(\u_fir|taps_13__15_ ),
	.datac(vcc),
	.datad(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hC33C;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N30
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|taps_14__15_  $ \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(\u_fir|taps_14__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hA55A;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N30
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  $ \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(vcc),
	.datab(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1 ),
	.datac(vcc),
	.datad(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hC33C;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N30
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|taps_16__15_  $ \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(\u_fir|taps_16__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hA55A;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N30
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52923 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z1  = \u_fir|tap_array_17_filter_block_tap_next_15_  $ \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z4  $ \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z1 

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z1 ),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z4 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52923 .lut_mask = 16'hA55A;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X33_Y2_N13
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_0_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx51271z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z17 ));

// atom is at LCFF_X33_Y2_N21
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_4_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx55259z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z9 ));

// atom is at LCFF_X33_Y2_N17
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_2_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx53265z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z13 ));

// atom is at LCCOMB_X34_Y2_N12
cycloneii_lcell_comb ix50205z52926(
// Equation(s):
// nx50205z4 = !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z7  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z9  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z11  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z13 

	.dataa(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z13 ),
	.datab(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z11 ),
	.datac(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z9 ),
	.datad(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z7 ),
	.cin(gnd),
	.combout(nx50205z4),
	.cout());
// synopsys translate_off
defparam ix50205z52926.lut_mask = 16'h7FFF;
defparam ix50205z52926.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X34_Y2_N6
cycloneii_lcell_comb ix50205z52925(
// Equation(s):
// nx50205z3 = nx50205z4 # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z17  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z15 

	.dataa(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z15 ),
	.datab(vcc),
	.datac(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z17 ),
	.datad(nx50205z4),
	.cin(gnd),
	.combout(nx50205z3),
	.cout());
// synopsys translate_off
defparam ix50205z52925.lut_mask = 16'hFF5F;
defparam ix50205z52925.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N13
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_4_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx55259z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z17 ));

// atom is at LCFF_X60_Y19_N29
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_12_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx1963z1 ));

// atom is at LCFF_X60_Y19_N17
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_6_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx57253z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z13 ));

// atom is at LCCOMB_X57_Y19_N18
cycloneii_lcell_comb \u_i2c_av_config|u0|ix44942z52930 (
// Equation(s):
// \u_i2c_av_config|u0|nx44942z8  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 

	.dataa(vcc),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx44942z8 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix44942z52930 .lut_mask = 16'h3F3F;
defparam \u_i2c_av_config|u0|ix44942z52930 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N10
cycloneii_lcell_comb \u_i2c_av_config|u0|ix7286z52924 (
// Equation(s):
// \u_i2c_av_config|u0|nx7286z2  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  # 
// !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx7286z2 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix7286z52924 .lut_mask = 16'h7FFF;
defparam \u_i2c_av_config|u0|ix7286z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X27_Y14_N7
cycloneii_lcell_ff u_sine_reg_address_0_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx37973z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_0_));

// atom is at LCCOMB_X27_Y14_N6
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52932 (
// Equation(s):
// \u_sine_address_add9_0i1|nx37973z1  = u_sine_address_0_ & (\sw~combout [0] # GND) # !u_sine_address_0_ & (\sw~combout [0] $ VCC)
// \u_sine_address_add9_0i1|nx45949z23  = CARRY(u_sine_address_0_ # \sw~combout [0])

	.dataa(u_sine_address_0_),
	.datab(\sw~combout [0]),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_sine_address_add9_0i1|nx37973z1 ),
	.cout(\u_sine_address_add9_0i1|nx45949z23 ));
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52932 .lut_mask = 16'h99EE;
defparam \u_sine_address_add9_0i1|ix45949z52932 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X27_Y14_N15
cycloneii_lcell_ff u_sine_reg_address_4_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx41961z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_4_));

// atom is at LCFF_X27_Y14_N17
cycloneii_lcell_ff u_sine_reg_address_5_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx42958z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_5_));

// atom is at LCFF_X27_Y14_N21
cycloneii_lcell_ff u_sine_reg_address_7_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx44952z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_7_));

// atom is at LCCOMB_X33_Y2_N12
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52932 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx51271z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z17  $ VCC
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z16  = CARRY(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z17 )

	.dataa(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z17 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx51271z1 ),
	.cout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z16 ));
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52932 .lut_mask = 16'h55AA;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52932 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X33_Y2_N16
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52930 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx53265z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z13  & (\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z14  $ GND) # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z13  & 
// !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z14  & VCC
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z12  = CARRY(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z13  & !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z14 )

	.dataa(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z13 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z14 ),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx53265z1 ),
	.cout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z12 ));
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52930 .lut_mask = 16'hA50A;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X33_Y2_N20
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52928 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx55259z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z9  & (\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z10  $ GND) # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z9  & 
// !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z10  & VCC
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z8  = CARRY(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z9  & !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z10 )

	.dataa(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z9 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z10 ),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx55259z1 ),
	.cout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z8 ));
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52928 .lut_mask = 16'hA50A;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N7
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_1_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx52268z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z23 ));

// atom is at LCCOMB_X60_Y19_N6
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52935 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx52268z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z23  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z24  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z23  & 
// (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z24  # GND)
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z22  = CARRY(!\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z24  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z23 )

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z23 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z24 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx52268z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z22 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52935 .lut_mask = 16'h5A5F;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y19_N12
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52932 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx55259z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z17  & (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z18  $ GND) # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z17  & 
// !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z18  & VCC
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z16  = CARRY(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z17  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z18 )

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z17 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z18 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx55259z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z16 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52932 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y19_N16
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52930 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx57253z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z13  & (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z14  $ GND) # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z13  & 
// !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z14  & VCC
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z12  = CARRY(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z13  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z14 )

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z13 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z14 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx57253z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z12 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52930 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y19_N26
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52925 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx18093z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z4  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3  & 
// (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z4  # GND)
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z2  = CARRY(!\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z4  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z4 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx18093z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z2 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52925 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y19_N28
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52923 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z2  $ !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx1963z1 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx1963z1 ),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z2 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52923 .lut_mask = 16'hF00F;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N11
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_5_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx56256z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_5_ ));

// atom is at LCFF_X54_Y19_N13
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_6_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx57253z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_6_ ));

// atom is at LCCOMB_X55_Y19_N6
cycloneii_lcell_comb \u_i2c_av_config|ix35560z52924 (
// Equation(s):
// \u_i2c_av_config|nx35560z2  = \u_i2c_av_config|modgen_counter_cont|q_6_  & \u_i2c_av_config|modgen_counter_cont|q_5_  & \u_i2c_av_config|modgen_counter_cont|q_7_  & \u_i2c_av_config|modgen_counter_cont|q_4_ 

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_6_ ),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_5_ ),
	.datac(\u_i2c_av_config|modgen_counter_cont|q_7_ ),
	.datad(\u_i2c_av_config|modgen_counter_cont|q_4_ ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx35560z2 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix35560z52924 .lut_mask = 16'h8000;
defparam \u_i2c_av_config|ix35560z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N24
cycloneii_lcell_comb \u_i2c_av_config|u0|ix22137z52926 (
// Equation(s):
// \u_i2c_av_config|u0|nx22137z2  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  & (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  # \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & 
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx22137z2 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix22137z52926 .lut_mask = 16'hF080;
defparam \u_i2c_av_config|u0|ix22137z52926 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N18
cycloneii_lcell_comb \u_i2c_av_config|u0|ix22137z52925 (
// Equation(s):
// \u_i2c_av_config|u0|sdo_5n5s2f1_0_  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  & (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  & !\u_i2c_av_config|u0|nx44942z5  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  & 
// (\u_i2c_av_config|u0|nx22137z2 ))

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datab(\u_i2c_av_config|u0|nx44942z5 ),
	.datac(\u_i2c_av_config|u0|nx22137z2 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|sdo_5n5s2f1_0_ ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix22137z52925 .lut_mask = 16'h1150;
defparam \u_i2c_av_config|u0|ix22137z52925 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N0
cycloneii_lcell_comb \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52928 (
// Equation(s):
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1  = \u_i2c_av_config|u0|sdo_5n5s2f1_0_  & (GND # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ) # !\u_i2c_av_config|u0|sdo_5n5s2f1_0_  & (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  $ 
// GND)
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11  = CARRY(\u_i2c_av_config|u0|sdo_5n5s2f1_0_  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 )

	.dataa(\u_i2c_av_config|u0|sdo_5n5s2f1_0_ ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1 ),
	.cout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52928 .lut_mask = 16'h66BB;
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52928 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N6
cycloneii_lcell_comb \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52925 (
// Equation(s):
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx40964z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z5  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  & \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z5  
// & VCC
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z3  = CARRY(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z5 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z5 ),
	.combout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx40964z1 ),
	.cout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z3 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52925 .lut_mask = 16'h5A0A;
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y19_N12
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52926 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z4  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  # !\u_i2c_av_config|u0|nx7286z2 

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datab(vcc),
	.datac(\u_i2c_av_config|u0|nx7286z2 ),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z4 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52926 .lut_mask = 16'hAFAF;
defparam \u_i2c_av_config|u0|ix41315z52926 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N10
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52932 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z10  = !\u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1  & (\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1  $ \u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1 ),
	.datac(\u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1 ),
	.datad(\u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z10 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52932 .lut_mask = 16'h030C;
defparam \u_i2c_av_config|u0|ix41315z52932 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N26
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52934 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z12  = !\u_i2c_av_config|u0|nx44942z4  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & !\u_i2c_av_config|u0|nx44942z7 

	.dataa(\u_i2c_av_config|u0|nx44942z4 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datad(\u_i2c_av_config|u0|nx44942z7 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z12 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52934 .lut_mask = 16'h0004;
defparam \u_i2c_av_config|u0|ix41315z52934 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N28
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52936 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z14  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 

	.dataa(vcc),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z14 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52936 .lut_mask = 16'h3000;
defparam \u_i2c_av_config|u0|ix41315z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N22
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52935 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z13  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & \u_i2c_av_config|u0|nx41315z14  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datab(\u_i2c_av_config|u0|nx41315z14 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z13 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52935 .lut_mask = 16'h0004;
defparam \u_i2c_av_config|u0|ix41315z52935 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N0
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52938 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z16  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datab(vcc),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z16 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52938 .lut_mask = 16'h0005;
defparam \u_i2c_av_config|u0|ix41315z52938 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N10
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52939 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z17  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & \u_i2c_av_config|u0|nx41315z14  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datab(\u_i2c_av_config|u0|nx41315z14 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z17 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52939 .lut_mask = 16'h4000;
defparam \u_i2c_av_config|u0|ix41315z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N20
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52937 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z15  = \u_i2c_av_config|u0|nx41315z17  # \u_i2c_av_config|u0|nx41315z16  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 

	.dataa(\u_i2c_av_config|u0|nx41315z17 ),
	.datab(\u_i2c_av_config|u0|nx41315z16 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z15 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52937 .lut_mask = 16'hAAAE;
defparam \u_i2c_av_config|u0|ix41315z52937 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N6
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52933 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z11  = \u_i2c_av_config|u0|nx41315z13  # \u_i2c_av_config|u0|nx41315z15  # \u_i2c_av_config|u0|nx41315z12 

	.dataa(vcc),
	.datab(\u_i2c_av_config|u0|nx41315z13 ),
	.datac(\u_i2c_av_config|u0|nx41315z15 ),
	.datad(\u_i2c_av_config|u0|nx41315z12 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z11 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52933 .lut_mask = 16'hFFFC;
defparam \u_i2c_av_config|u0|ix41315z52933 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N16
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52943 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z21  = !\u_i2c_av_config|u0|nx44942z4  & !\u_i2c_av_config|u0|nx44942z5  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 

	.dataa(\u_i2c_av_config|u0|nx44942z4 ),
	.datab(\u_i2c_av_config|u0|nx44942z5 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z21 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52943 .lut_mask = 16'h0100;
defparam \u_i2c_av_config|u0|ix41315z52943 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N2
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52944 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z22  = \u_i2c_av_config|u0|nx41315z15  # !\u_i2c_av_config|u0|nx44942z7  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & \u_i2c_av_config|u0|nx41315z14 

	.dataa(\u_i2c_av_config|u0|nx41315z15 ),
	.datab(\u_i2c_av_config|u0|nx44942z7 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datad(\u_i2c_av_config|u0|nx41315z14 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z22 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52944 .lut_mask = 16'hABAA;
defparam \u_i2c_av_config|u0|ix41315z52944 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N12
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52942 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z20  = !\u_i2c_av_config|u0|nx41315z21  & (\u_i2c_av_config|u0|nx41315z22  # !\u_i2c_av_config|u0|nx41315z4 ) # !\u_i2c_av_config|reset_n 

	.dataa(\u_i2c_av_config|reset_n ),
	.datab(\u_i2c_av_config|u0|nx41315z22 ),
	.datac(\u_i2c_av_config|u0|nx41315z21 ),
	.datad(\u_i2c_av_config|u0|nx41315z4 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z20 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52942 .lut_mask = 16'h5D5F;
defparam \u_i2c_av_config|u0|ix41315z52942 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X54_Y19_N10
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52934 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx56256z1  = \u_i2c_av_config|modgen_counter_cont|q_5_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z12  # !\u_i2c_av_config|modgen_counter_cont|q_5_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z12  # GND)
// \u_i2c_av_config|modgen_counter_cont|nx22081z11  = CARRY(!\u_i2c_av_config|modgen_counter_cont|nx22081z12  # !\u_i2c_av_config|modgen_counter_cont|q_5_ )

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_5_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z12 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx56256z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z11 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52934 .lut_mask = 16'h5A5F;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y19_N12
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52933 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx57253z1  = \u_i2c_av_config|modgen_counter_cont|q_6_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z11  $ GND) # !\u_i2c_av_config|modgen_counter_cont|q_6_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z11  & VCC
// \u_i2c_av_config|modgen_counter_cont|nx22081z10  = CARRY(\u_i2c_av_config|modgen_counter_cont|q_6_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z11 )

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_6_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z11 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx57253z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z10 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52933 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at CLKCTRL_G15
cycloneii_clkctrl \aud_bclk_dup0~clkctrl (
	.ena(vcc),
	.inclk({gnd,gnd,gnd,aud_bclk_dup0}),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\aud_bclk_dup0~clkctrl_outclk ));
// synopsys translate_off
defparam \aud_bclk_dup0~clkctrl .clock_type = "global clock";
defparam \aud_bclk_dup0~clkctrl .ena_register_mode = "falling edge";
// synopsys translate_on

// atom is at LCCOMB_X34_Y14_N6
cycloneii_lcell_comb \audio_out_0_~feeder (
// Equation(s):
// \audio_out_0_~feeder_combout  = raw_audio_0_

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(raw_audio_0_),
	.cin(gnd),
	.combout(\audio_out_0_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \audio_out_0_~feeder .lut_mask = 16'hFF00;
defparam \audio_out_0_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X35_Y14_N10
cycloneii_lcell_comb \audio_out_15_~feeder (
// Equation(s):
// \audio_out_15_~feeder_combout  = raw_audio_11_

	.dataa(vcc),
	.datab(raw_audio_11_),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\audio_out_15_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \audio_out_15_~feeder .lut_mask = 16'hCCCC;
defparam \audio_out_15_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at PIN_N25
cycloneii_io sw_ibuf_0_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [0]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[0]));
// synopsys translate_off
defparam sw_ibuf_0_.input_async_reset = "none";
defparam sw_ibuf_0_.input_power_up = "low";
defparam sw_ibuf_0_.input_register_mode = "none";
defparam sw_ibuf_0_.input_sync_reset = "none";
defparam sw_ibuf_0_.oe_async_reset = "none";
defparam sw_ibuf_0_.oe_power_up = "low";
defparam sw_ibuf_0_.oe_register_mode = "none";
defparam sw_ibuf_0_.oe_sync_reset = "none";
defparam sw_ibuf_0_.operation_mode = "input";
defparam sw_ibuf_0_.output_async_reset = "none";
defparam sw_ibuf_0_.output_power_up = "low";
defparam sw_ibuf_0_.output_register_mode = "none";
defparam sw_ibuf_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AE14
cycloneii_io sw_ibuf_3_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [3]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[3]));
// synopsys translate_off
defparam sw_ibuf_3_.input_async_reset = "none";
defparam sw_ibuf_3_.input_power_up = "low";
defparam sw_ibuf_3_.input_register_mode = "none";
defparam sw_ibuf_3_.input_sync_reset = "none";
defparam sw_ibuf_3_.oe_async_reset = "none";
defparam sw_ibuf_3_.oe_power_up = "low";
defparam sw_ibuf_3_.oe_register_mode = "none";
defparam sw_ibuf_3_.oe_sync_reset = "none";
defparam sw_ibuf_3_.operation_mode = "input";
defparam sw_ibuf_3_.output_async_reset = "none";
defparam sw_ibuf_3_.output_power_up = "low";
defparam sw_ibuf_3_.output_register_mode = "none";
defparam sw_ibuf_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P25
cycloneii_io sw_ibuf_2_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [2]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[2]));
// synopsys translate_off
defparam sw_ibuf_2_.input_async_reset = "none";
defparam sw_ibuf_2_.input_power_up = "low";
defparam sw_ibuf_2_.input_register_mode = "none";
defparam sw_ibuf_2_.input_sync_reset = "none";
defparam sw_ibuf_2_.oe_async_reset = "none";
defparam sw_ibuf_2_.oe_power_up = "low";
defparam sw_ibuf_2_.oe_register_mode = "none";
defparam sw_ibuf_2_.oe_sync_reset = "none";
defparam sw_ibuf_2_.operation_mode = "input";
defparam sw_ibuf_2_.output_async_reset = "none";
defparam sw_ibuf_2_.output_power_up = "low";
defparam sw_ibuf_2_.output_register_mode = "none";
defparam sw_ibuf_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N30
cycloneii_lcell_comb ix49625z52929(
// Equation(s):
// nx49625z3 = \sw~combout [1] & !\sw~combout [2] & (\sw~combout [0] # \sw~combout [3]) # !\sw~combout [1] & (\sw~combout [3] & \sw~combout [0] & !\sw~combout [2] # !\sw~combout [3] & (\sw~combout [2]))

	.dataa(\sw~combout [1]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx49625z3),
	.cout());
// synopsys translate_off
defparam ix49625z52929.lut_mask = 16'h05E8;
defparam ix49625z52929.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at PIN_V2
cycloneii_io sw_ibuf_17_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [17]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[17]));
// synopsys translate_off
defparam sw_ibuf_17_.input_async_reset = "none";
defparam sw_ibuf_17_.input_power_up = "low";
defparam sw_ibuf_17_.input_register_mode = "none";
defparam sw_ibuf_17_.input_sync_reset = "none";
defparam sw_ibuf_17_.oe_async_reset = "none";
defparam sw_ibuf_17_.oe_power_up = "low";
defparam sw_ibuf_17_.oe_register_mode = "none";
defparam sw_ibuf_17_.oe_sync_reset = "none";
defparam sw_ibuf_17_.operation_mode = "input";
defparam sw_ibuf_17_.output_async_reset = "none";
defparam sw_ibuf_17_.output_power_up = "low";
defparam sw_ibuf_17_.output_register_mode = "none";
defparam sw_ibuf_17_.output_sync_reset = "none";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N12
cycloneii_lcell_comb ix49625z52925(
// Equation(s):
// nx49625z1 = \sw~combout [3] & \sw~combout [1] & \sw~combout [0] & \sw~combout [2] # !\sw~combout [3] & !\sw~combout [2] & (!\sw~combout [0] # !\sw~combout [1])

	.dataa(\sw~combout [1]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx49625z1),
	.cout());
// synopsys translate_off
defparam ix49625z52925.lut_mask = 16'h8007;
defparam ix49625z52925.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X34_Y14_N26
cycloneii_lcell_comb ix55607z52924(
// Equation(s):
// nx55607z1 = nx49625z2 & !nx49625z3 & !\sw~combout [17] & !nx49625z1

	.dataa(nx49625z2),
	.datab(nx49625z3),
	.datac(\sw~combout [17]),
	.datad(nx49625z1),
	.cin(gnd),
	.combout(nx55607z1),
	.cout());
// synopsys translate_off
defparam ix55607z52924.lut_mask = 16'h0002;
defparam ix55607z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N2
cycloneii_lcell_comb ix49625z52931(
// Equation(s):
// nx49625z4 = \sw~combout [3] $ (\sw~combout [1] & (\sw~combout [0] $ \sw~combout [2]) # !\sw~combout [1] & !\sw~combout [0] & !\sw~combout [2])

	.dataa(\sw~combout [1]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx49625z4),
	.cout());
// synopsys translate_off
defparam ix49625z52931.lut_mask = 16'hD269;
defparam ix49625z52931.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X34_Y14_N24
cycloneii_lcell_comb ix49625z52930(
// Equation(s):
// display_freq_0_ = !\sw~combout [17] & nx49625z4

	.dataa(vcc),
	.datab(vcc),
	.datac(\sw~combout [17]),
	.datad(nx49625z4),
	.cin(gnd),
	.combout(display_freq_0_),
	.cout());
// synopsys translate_off
defparam ix49625z52930.lut_mask = 16'h0F00;
defparam ix49625z52930.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N24
cycloneii_lcell_comb ix49625z52928(
// Equation(s):
// display_freq_1_ = \sw~combout [17] # nx49625z3

	.dataa(vcc),
	.datab(\sw~combout [17]),
	.datac(vcc),
	.datad(nx49625z3),
	.cin(gnd),
	.combout(display_freq_1_),
	.cout());
// synopsys translate_off
defparam ix49625z52928.lut_mask = 16'hFFCC;
defparam ix49625z52928.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N8
cycloneii_lcell_comb ix49625z52927(
// Equation(s):
// nx49625z2 = \sw~combout [3] & !\sw~combout [1] & !\sw~combout [0] & !\sw~combout [2] # !\sw~combout [3] & (\sw~combout [2] # \sw~combout [1] & \sw~combout [0])

	.dataa(\sw~combout [1]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx49625z2),
	.cout());
// synopsys translate_off
defparam ix49625z52927.lut_mask = 16'h0F18;
defparam ix49625z52927.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N26
cycloneii_lcell_comb ix49625z52926(
// Equation(s):
// display_freq_2_ = \sw~combout [17] # nx49625z2

	.dataa(\sw~combout [17]),
	.datab(vcc),
	.datac(vcc),
	.datad(nx49625z2),
	.cin(gnd),
	.combout(display_freq_2_),
	.cout());
// synopsys translate_off
defparam ix49625z52926.lut_mask = 16'hFFAA;
defparam ix49625z52926.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y14_N0
cycloneii_lcell_comb ix55607z52925(
// Equation(s):
// nx55607z2 = display_freq_0_ & (display_freq_3_ & (display_freq_1_ $ display_freq_2_) # !display_freq_3_ & !display_freq_1_ & !display_freq_2_)

	.dataa(display_freq_3_),
	.datab(display_freq_0_),
	.datac(display_freq_1_),
	.datad(display_freq_2_),
	.cin(gnd),
	.combout(nx55607z2),
	.cout());
// synopsys translate_off
defparam ix55607z52925.lut_mask = 16'h0884;
defparam ix55607z52925.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y14_N18
cycloneii_lcell_comb ix55607z52923(
// Equation(s):
// hex4_dup0_0_ = nx55607z2 # nx55607z1 & !display_freq_0_ & display_freq_2_

	.dataa(nx55607z1),
	.datab(nx55607z2),
	.datac(display_freq_0_),
	.datad(display_freq_2_),
	.cin(gnd),
	.combout(hex4_dup0_0_),
	.cout());
// synopsys translate_off
defparam ix55607z52923.lut_mask = 16'hCECC;
defparam ix55607z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X34_Y14_N20
cycloneii_lcell_comb ix49625z52924(
// Equation(s):
// display_freq_3_ = \sw~combout [17] # nx49625z1

	.dataa(vcc),
	.datab(vcc),
	.datac(\sw~combout [17]),
	.datad(nx49625z1),
	.cin(gnd),
	.combout(display_freq_3_),
	.cout());
// synopsys translate_off
defparam ix49625z52924.lut_mask = 16'hFFF0;
defparam ix49625z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y14_N20
cycloneii_lcell_comb ix54610z52923(
// Equation(s):
// hex4_dup0_1_ = display_freq_3_ & (display_freq_0_ & display_freq_1_ # !display_freq_0_ & (display_freq_2_)) # !display_freq_3_ & display_freq_2_ & (display_freq_0_ $ display_freq_1_)

	.dataa(display_freq_3_),
	.datab(display_freq_0_),
	.datac(display_freq_1_),
	.datad(display_freq_2_),
	.cin(gnd),
	.combout(hex4_dup0_1_),
	.cout());
// synopsys translate_off
defparam ix54610z52923.lut_mask = 16'hB680;
defparam ix54610z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y14_N22
cycloneii_lcell_comb ix53613z52923(
// Equation(s):
// hex4_dup0_2_ = display_freq_3_ & display_freq_2_ & (display_freq_1_ # !display_freq_0_) # !display_freq_3_ & !display_freq_0_ & display_freq_1_ & !display_freq_2_

	.dataa(display_freq_3_),
	.datab(display_freq_0_),
	.datac(display_freq_1_),
	.datad(display_freq_2_),
	.cin(gnd),
	.combout(hex4_dup0_2_),
	.cout());
// synopsys translate_off
defparam ix53613z52923.lut_mask = 16'hA210;
defparam ix53613z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y14_N24
cycloneii_lcell_comb ix52616z52923(
// Equation(s):
// hex4_dup0_3_ = display_freq_0_ & (display_freq_1_ $ !display_freq_2_) # !display_freq_0_ & (display_freq_3_ & display_freq_1_ & !display_freq_2_ # !display_freq_3_ & !display_freq_1_ & display_freq_2_)

	.dataa(display_freq_3_),
	.datab(display_freq_0_),
	.datac(display_freq_1_),
	.datad(display_freq_2_),
	.cin(gnd),
	.combout(hex4_dup0_3_),
	.cout());
// synopsys translate_off
defparam ix52616z52923.lut_mask = 16'hC12C;
defparam ix52616z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y14_N26
cycloneii_lcell_comb ix51619z52923(
// Equation(s):
// hex4_dup0_4_ = display_freq_1_ & !display_freq_3_ & display_freq_0_ # !display_freq_1_ & (display_freq_2_ & !display_freq_3_ # !display_freq_2_ & (display_freq_0_))

	.dataa(display_freq_3_),
	.datab(display_freq_0_),
	.datac(display_freq_1_),
	.datad(display_freq_2_),
	.cin(gnd),
	.combout(hex4_dup0_4_),
	.cout());
// synopsys translate_off
defparam ix51619z52923.lut_mask = 16'h454C;
defparam ix51619z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y14_N28
cycloneii_lcell_comb ix50622z52923(
// Equation(s):
// hex4_dup0_5_ = display_freq_0_ & (display_freq_3_ $ (display_freq_1_ # !display_freq_2_)) # !display_freq_0_ & !display_freq_3_ & display_freq_1_ & !display_freq_2_

	.dataa(display_freq_3_),
	.datab(display_freq_0_),
	.datac(display_freq_1_),
	.datad(display_freq_2_),
	.cin(gnd),
	.combout(hex4_dup0_5_),
	.cout());
// synopsys translate_off
defparam ix50622z52923.lut_mask = 16'h4854;
defparam ix50622z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y14_N6
cycloneii_lcell_comb ix49625z52923(
// Equation(s):
// hex4_dup0_6_ = display_freq_0_ & !display_freq_3_ & (display_freq_1_ $ !display_freq_2_) # !display_freq_0_ & !display_freq_1_ & (display_freq_3_ $ !display_freq_2_)

	.dataa(display_freq_3_),
	.datab(display_freq_0_),
	.datac(display_freq_1_),
	.datad(display_freq_2_),
	.cin(gnd),
	.combout(hex4_dup0_6_),
	.cout());
// synopsys translate_off
defparam ix49625z52923.lut_mask = 16'h4205;
defparam ix49625z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at PIN_AF14
cycloneii_io sw_ibuf_4_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [4]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[4]));
// synopsys translate_off
defparam sw_ibuf_4_.input_async_reset = "none";
defparam sw_ibuf_4_.input_power_up = "low";
defparam sw_ibuf_4_.input_register_mode = "none";
defparam sw_ibuf_4_.input_sync_reset = "none";
defparam sw_ibuf_4_.oe_async_reset = "none";
defparam sw_ibuf_4_.oe_power_up = "low";
defparam sw_ibuf_4_.oe_register_mode = "none";
defparam sw_ibuf_4_.oe_sync_reset = "none";
defparam sw_ibuf_4_.operation_mode = "input";
defparam sw_ibuf_4_.output_async_reset = "none";
defparam sw_ibuf_4_.output_power_up = "low";
defparam sw_ibuf_4_.output_register_mode = "none";
defparam sw_ibuf_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_N26
cycloneii_io sw_ibuf_1_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [1]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[1]));
// synopsys translate_off
defparam sw_ibuf_1_.input_async_reset = "none";
defparam sw_ibuf_1_.input_power_up = "low";
defparam sw_ibuf_1_.input_register_mode = "none";
defparam sw_ibuf_1_.input_sync_reset = "none";
defparam sw_ibuf_1_.oe_async_reset = "none";
defparam sw_ibuf_1_.oe_power_up = "low";
defparam sw_ibuf_1_.oe_register_mode = "none";
defparam sw_ibuf_1_.oe_sync_reset = "none";
defparam sw_ibuf_1_.operation_mode = "input";
defparam sw_ibuf_1_.output_async_reset = "none";
defparam sw_ibuf_1_.output_power_up = "low";
defparam sw_ibuf_1_.output_register_mode = "none";
defparam sw_ibuf_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N18
cycloneii_lcell_comb ix38664z52935(
// Equation(s):
// nx38664z8 = \sw~combout [3] & (\sw~combout [1] & nx38664z9 # !\sw~combout [1] & (\sw~combout [4])) # !\sw~combout [3] & (\sw~combout [4])

	.dataa(nx38664z9),
	.datab(\sw~combout [4]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [1]),
	.cin(gnd),
	.combout(nx38664z8),
	.cout());
// synopsys translate_off
defparam ix38664z52935.lut_mask = 16'hACCC;
defparam ix38664z52935.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N12
cycloneii_lcell_comb ix38664z52934(
// Equation(s):
// display_freq_4_ = \sw~combout [17] # \sw~combout [0] & nx38664z8 # !\sw~combout [0] & (!\sw~combout [4])

	.dataa(\sw~combout [17]),
	.datab(nx38664z8),
	.datac(\sw~combout [4]),
	.datad(\sw~combout [0]),
	.cin(gnd),
	.combout(display_freq_4_),
	.cout());
// synopsys translate_off
defparam ix38664z52934.lut_mask = 16'hEEAF;
defparam ix38664z52934.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N20
cycloneii_lcell_comb ix38664z52926(
// Equation(s):
// nx38664z2 = \sw~combout [3] & !\sw~combout [0] & !\sw~combout [1] & !\sw~combout [4] # !\sw~combout [3] & (\sw~combout [1] & \sw~combout [4])

	.dataa(\sw~combout [3]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [1]),
	.datad(\sw~combout [4]),
	.cin(gnd),
	.combout(nx38664z2),
	.cout());
// synopsys translate_off
defparam ix38664z52926.lut_mask = 16'h5002;
defparam ix38664z52926.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N6
cycloneii_lcell_comb ix38664z52924(
// Equation(s):
// display_freq_7_ = !\sw~combout [17] & (\sw~combout [2] & nx38664z1 # !\sw~combout [2] & (nx38664z2))

	.dataa(nx38664z1),
	.datab(\sw~combout [17]),
	.datac(nx38664z2),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(display_freq_7_),
	.cout());
// synopsys translate_off
defparam ix38664z52924.lut_mask = 16'h2230;
defparam ix38664z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at PIN_AC13
cycloneii_io sw_ibuf_6_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [6]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[6]));
// synopsys translate_off
defparam sw_ibuf_6_.input_async_reset = "none";
defparam sw_ibuf_6_.input_power_up = "low";
defparam sw_ibuf_6_.input_register_mode = "none";
defparam sw_ibuf_6_.input_sync_reset = "none";
defparam sw_ibuf_6_.oe_async_reset = "none";
defparam sw_ibuf_6_.oe_power_up = "low";
defparam sw_ibuf_6_.oe_register_mode = "none";
defparam sw_ibuf_6_.oe_sync_reset = "none";
defparam sw_ibuf_6_.operation_mode = "input";
defparam sw_ibuf_6_.output_async_reset = "none";
defparam sw_ibuf_6_.output_power_up = "low";
defparam sw_ibuf_6_.output_register_mode = "none";
defparam sw_ibuf_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N24
cycloneii_lcell_comb ix38664z52930(
// Equation(s):
// nx38664z5 = !\sw~combout [2] & (\sw~combout [5] # !\sw~combout [6] # !\sw~combout [0])

	.dataa(\sw~combout [5]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [6]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx38664z5),
	.cout());
// synopsys translate_off
defparam ix38664z52930.lut_mask = 16'h00BF;
defparam ix38664z52930.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N26
cycloneii_lcell_comb ix38664z52929(
// Equation(s):
// nx38664z4 = \sw~combout [1] & \sw~combout [3] & nx38664z5 # !\sw~combout [1] & (!\sw~combout [2])

	.dataa(\sw~combout [3]),
	.datab(nx38664z5),
	.datac(\sw~combout [1]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx38664z4),
	.cout());
// synopsys translate_off
defparam ix38664z52929.lut_mask = 16'h808F;
defparam ix38664z52929.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N0
cycloneii_lcell_comb ix38664z52927(
// Equation(s):
// display_freq_6_ = \sw~combout [17] # \sw~combout [4] & (nx38664z4) # !\sw~combout [4] & nx38664z3

	.dataa(nx38664z3),
	.datab(nx38664z4),
	.datac(\sw~combout [4]),
	.datad(\sw~combout [17]),
	.cin(gnd),
	.combout(display_freq_6_),
	.cout());
// synopsys translate_off
defparam ix38664z52927.lut_mask = 16'hFFCA;
defparam ix38664z52927.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N4
cycloneii_lcell_comb ix38664z52932(
// Equation(s):
// nx38664z6 = \sw~combout [3] & !\sw~combout [0] & !\sw~combout [1] & !\sw~combout [4] # !\sw~combout [3] & (\sw~combout [1] $ (\sw~combout [0] & !\sw~combout [4]))

	.dataa(\sw~combout [3]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [1]),
	.datad(\sw~combout [4]),
	.cin(gnd),
	.combout(nx38664z6),
	.cout());
// synopsys translate_off
defparam ix38664z52932.lut_mask = 16'h5016;
defparam ix38664z52932.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N14
cycloneii_lcell_comb ix38664z52933(
// Equation(s):
// nx38664z7 = \sw~combout [3] & \sw~combout [1] & (\sw~combout [0] # \sw~combout [4]) # !\sw~combout [3] & (\sw~combout [1] $ (\sw~combout [0] # \sw~combout [4]))

	.dataa(\sw~combout [3]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [1]),
	.datad(\sw~combout [4]),
	.cin(gnd),
	.combout(nx38664z7),
	.cout());
// synopsys translate_off
defparam ix38664z52933.lut_mask = 16'hA594;
defparam ix38664z52933.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N0
cycloneii_lcell_comb ix38664z52931(
// Equation(s):
// display_freq_5_ = !\sw~combout [17] & (\sw~combout [2] & nx38664z6 # !\sw~combout [2] & (nx38664z7))

	.dataa(\sw~combout [17]),
	.datab(nx38664z6),
	.datac(nx38664z7),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(display_freq_5_),
	.cout());
// synopsys translate_off
defparam ix38664z52931.lut_mask = 16'h4450;
defparam ix38664z52931.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y15_N24
cycloneii_lcell_comb ix32682z52923(
// Equation(s):
// hex5_dup0_0_ = display_freq_7_ & display_freq_4_ & (display_freq_6_ $ display_freq_5_) # !display_freq_7_ & !display_freq_5_ & (display_freq_4_ $ display_freq_6_)

	.dataa(display_freq_4_),
	.datab(display_freq_7_),
	.datac(display_freq_6_),
	.datad(display_freq_5_),
	.cin(gnd),
	.combout(hex5_dup0_0_),
	.cout());
// synopsys translate_off
defparam ix32682z52923.lut_mask = 16'h0892;
defparam ix32682z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y15_N26
cycloneii_lcell_comb ix33679z52923(
// Equation(s):
// hex5_dup0_1_ = display_freq_7_ & (display_freq_4_ & (display_freq_5_) # !display_freq_4_ & display_freq_6_) # !display_freq_7_ & display_freq_6_ & (display_freq_4_ $ display_freq_5_)

	.dataa(display_freq_4_),
	.datab(display_freq_7_),
	.datac(display_freq_6_),
	.datad(display_freq_5_),
	.cin(gnd),
	.combout(hex5_dup0_1_),
	.cout());
// synopsys translate_off
defparam ix33679z52923.lut_mask = 16'hD860;
defparam ix33679z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y15_N20
cycloneii_lcell_comb ix34676z52923(
// Equation(s):
// hex5_dup0_2_ = display_freq_7_ & display_freq_6_ & (display_freq_5_ # !display_freq_4_) # !display_freq_7_ & !display_freq_4_ & !display_freq_6_ & display_freq_5_

	.dataa(display_freq_4_),
	.datab(display_freq_7_),
	.datac(display_freq_6_),
	.datad(display_freq_5_),
	.cin(gnd),
	.combout(hex5_dup0_2_),
	.cout());
// synopsys translate_off
defparam ix34676z52923.lut_mask = 16'hC140;
defparam ix34676z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y15_N22
cycloneii_lcell_comb ix35673z52923(
// Equation(s):
// hex5_dup0_3_ = display_freq_4_ & (display_freq_6_ $ !display_freq_5_) # !display_freq_4_ & (display_freq_7_ & !display_freq_6_ & display_freq_5_ # !display_freq_7_ & display_freq_6_ & !display_freq_5_)

	.dataa(display_freq_4_),
	.datab(display_freq_7_),
	.datac(display_freq_6_),
	.datad(display_freq_5_),
	.cin(gnd),
	.combout(hex5_dup0_3_),
	.cout());
// synopsys translate_off
defparam ix35673z52923.lut_mask = 16'hA41A;
defparam ix35673z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y15_N0
cycloneii_lcell_comb ix36670z52923(
// Equation(s):
// hex5_dup0_4_ = display_freq_5_ & display_freq_4_ & !display_freq_7_ # !display_freq_5_ & (display_freq_6_ & (!display_freq_7_) # !display_freq_6_ & display_freq_4_)

	.dataa(display_freq_4_),
	.datab(display_freq_7_),
	.datac(display_freq_6_),
	.datad(display_freq_5_),
	.cin(gnd),
	.combout(hex5_dup0_4_),
	.cout());
// synopsys translate_off
defparam ix36670z52923.lut_mask = 16'h223A;
defparam ix36670z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y15_N10
cycloneii_lcell_comb ix37667z52923(
// Equation(s):
// hex5_dup0_5_ = display_freq_4_ & (display_freq_7_ $ (display_freq_5_ # !display_freq_6_)) # !display_freq_4_ & !display_freq_7_ & !display_freq_6_ & display_freq_5_

	.dataa(display_freq_4_),
	.datab(display_freq_7_),
	.datac(display_freq_6_),
	.datad(display_freq_5_),
	.cin(gnd),
	.combout(hex5_dup0_5_),
	.cout());
// synopsys translate_off
defparam ix37667z52923.lut_mask = 16'h2382;
defparam ix37667z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y15_N12
cycloneii_lcell_comb ix38664z52923(
// Equation(s):
// hex5_dup0_6_ = display_freq_4_ & !display_freq_7_ & (display_freq_6_ $ !display_freq_5_) # !display_freq_4_ & !display_freq_5_ & (display_freq_7_ $ !display_freq_6_)

	.dataa(display_freq_4_),
	.datab(display_freq_7_),
	.datac(display_freq_6_),
	.datad(display_freq_5_),
	.cin(gnd),
	.combout(hex5_dup0_6_),
	.cout());
// synopsys translate_off
defparam ix38664z52923.lut_mask = 16'h2043;
defparam ix38664z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at PIN_AD13
cycloneii_io sw_ibuf_5_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [5]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[5]));
// synopsys translate_off
defparam sw_ibuf_5_.input_async_reset = "none";
defparam sw_ibuf_5_.input_power_up = "low";
defparam sw_ibuf_5_.input_register_mode = "none";
defparam sw_ibuf_5_.input_sync_reset = "none";
defparam sw_ibuf_5_.oe_async_reset = "none";
defparam sw_ibuf_5_.oe_power_up = "low";
defparam sw_ibuf_5_.oe_register_mode = "none";
defparam sw_ibuf_5_.oe_sync_reset = "none";
defparam sw_ibuf_5_.operation_mode = "input";
defparam sw_ibuf_5_.output_async_reset = "none";
defparam sw_ibuf_5_.output_power_up = "low";
defparam sw_ibuf_5_.output_register_mode = "none";
defparam sw_ibuf_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N18
cycloneii_lcell_comb ix4119z52932(
// Equation(s):
// nx4119z7 = \sw~combout [3] & (\sw~combout [1] # \sw~combout [0] # \sw~combout [2])

	.dataa(\sw~combout [1]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx4119z7),
	.cout());
// synopsys translate_off
defparam ix4119z52932.lut_mask = 16'hF0E0;
defparam ix4119z52932.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N16
cycloneii_lcell_comb ix4119z52931(
// Equation(s):
// nx4119z6 = \sw~combout [6] # \sw~combout [5] & (\sw~combout [4] # nx4119z7)

	.dataa(\sw~combout [6]),
	.datab(\sw~combout [4]),
	.datac(\sw~combout [5]),
	.datad(nx4119z7),
	.cin(gnd),
	.combout(nx4119z6),
	.cout());
// synopsys translate_off
defparam ix4119z52931.lut_mask = 16'hFAEA;
defparam ix4119z52931.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N30
cycloneii_lcell_comb ix4119z52930(
// Equation(s):
// nx4119z5 = !\sw~combout [5] & (!\sw~combout [3] & !\sw~combout [2] # !\sw~combout [4])

	.dataa(\sw~combout [5]),
	.datab(\sw~combout [4]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx4119z5),
	.cout());
// synopsys translate_off
defparam ix4119z52930.lut_mask = 16'h1115;
defparam ix4119z52930.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N26
cycloneii_lcell_comb ix4119z52929(
// Equation(s):
// display_freq_10_ = !\sw~combout [17] & nx4119z6 & (nx4119z5 # !\sw~combout [6])

	.dataa(\sw~combout [6]),
	.datab(\sw~combout [17]),
	.datac(nx4119z6),
	.datad(nx4119z5),
	.cin(gnd),
	.combout(display_freq_10_),
	.cout());
// synopsys translate_off
defparam ix4119z52929.lut_mask = 16'h3010;
defparam ix4119z52929.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N2
cycloneii_lcell_comb ix4119z52941(
// Equation(s):
// nx4119z14 = \sw~combout [4] # \sw~combout [3] & nx4119z15 # !\sw~combout [3] & (\sw~combout [5])

	.dataa(nx4119z15),
	.datab(\sw~combout [3]),
	.datac(\sw~combout [4]),
	.datad(\sw~combout [5]),
	.cin(gnd),
	.combout(nx4119z14),
	.cout());
// synopsys translate_off
defparam ix4119z52941.lut_mask = 16'hFBF8;
defparam ix4119z52941.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N20
cycloneii_lcell_comb ix4119z52939(
// Equation(s):
// display_freq_8_ = \sw~combout [17] # nx4119z14 & (nx4119z13 # !\sw~combout [4])

	.dataa(nx4119z13),
	.datab(\sw~combout [17]),
	.datac(\sw~combout [4]),
	.datad(nx4119z14),
	.cin(gnd),
	.combout(display_freq_8_),
	.cout());
// synopsys translate_off
defparam ix4119z52939.lut_mask = 16'hEFCC;
defparam ix4119z52939.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N28
cycloneii_lcell_comb ix4119z52934(
// Equation(s):
// nx4119z8 = \sw~combout [5] & !\sw~combout [6] & !\sw~combout [4] # !\sw~combout [5] & (\sw~combout [6] $ (\sw~combout [4] & \sw~combout [2]))

	.dataa(\sw~combout [5]),
	.datab(\sw~combout [6]),
	.datac(\sw~combout [4]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx4119z8),
	.cout());
// synopsys translate_off
defparam ix4119z52934.lut_mask = 16'h1646;
defparam ix4119z52934.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N4
cycloneii_lcell_comb ix4119z52933(
// Equation(s):
// display_freq_9_ = !\sw~combout [17] & (\sw~combout [3] & nx4119z9 # !\sw~combout [3] & (nx4119z8))

	.dataa(nx4119z9),
	.datab(nx4119z8),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [17]),
	.cin(gnd),
	.combout(display_freq_9_),
	.cout());
// synopsys translate_off
defparam ix4119z52933.lut_mask = 16'h00AC;
defparam ix4119z52933.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N14
cycloneii_lcell_comb ix4119z52925(
// Equation(s):
// nx4119z1 = \sw~combout [5] & !\sw~combout [4] # !\sw~combout [5] & \sw~combout [4] & \sw~combout [2]

	.dataa(vcc),
	.datab(\sw~combout [5]),
	.datac(\sw~combout [4]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx4119z1),
	.cout());
// synopsys translate_off
defparam ix4119z52925.lut_mask = 16'h3C0C;
defparam ix4119z52925.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X29_Y15_N8
cycloneii_lcell_comb ix4119z52928(
// Equation(s):
// nx4119z4 = \sw~combout [6] & !\sw~combout [17]

	.dataa(vcc),
	.datab(\sw~combout [6]),
	.datac(\sw~combout [17]),
	.datad(vcc),
	.cin(gnd),
	.combout(nx4119z4),
	.cout());
// synopsys translate_off
defparam ix4119z52928.lut_mask = 16'h0C0C;
defparam ix4119z52928.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N28
cycloneii_lcell_comb ix4119z52924(
// Equation(s):
// display_freq_11_ = nx4119z4 & (\sw~combout [3] & nx4119z2 # !\sw~combout [3] & (nx4119z1))

	.dataa(nx4119z2),
	.datab(nx4119z1),
	.datac(\sw~combout [3]),
	.datad(nx4119z4),
	.cin(gnd),
	.combout(display_freq_11_),
	.cout());
// synopsys translate_off
defparam ix4119z52924.lut_mask = 16'hAC00;
defparam ix4119z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y23_N24
cycloneii_lcell_comb ix10101z52923(
// Equation(s):
// hex6_dup0_0_ = display_freq_10_ & !display_freq_9_ & (display_freq_8_ $ !display_freq_11_) # !display_freq_10_ & display_freq_8_ & (display_freq_9_ $ !display_freq_11_)

	.dataa(display_freq_10_),
	.datab(display_freq_8_),
	.datac(display_freq_9_),
	.datad(display_freq_11_),
	.cin(gnd),
	.combout(hex6_dup0_0_),
	.cout());
// synopsys translate_off
defparam ix10101z52923.lut_mask = 16'h4806;
defparam ix10101z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y23_N10
cycloneii_lcell_comb ix9104z52923(
// Equation(s):
// hex6_dup0_1_ = display_freq_9_ & (display_freq_8_ & (display_freq_11_) # !display_freq_8_ & display_freq_10_) # !display_freq_9_ & display_freq_10_ & (display_freq_8_ $ display_freq_11_)

	.dataa(display_freq_10_),
	.datab(display_freq_8_),
	.datac(display_freq_9_),
	.datad(display_freq_11_),
	.cin(gnd),
	.combout(hex6_dup0_1_),
	.cout());
// synopsys translate_off
defparam ix9104z52923.lut_mask = 16'hE228;
defparam ix9104z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y23_N28
cycloneii_lcell_comb ix8107z52923(
// Equation(s):
// hex6_dup0_2_ = display_freq_10_ & display_freq_11_ & (display_freq_9_ # !display_freq_8_) # !display_freq_10_ & !display_freq_8_ & display_freq_9_ & !display_freq_11_

	.dataa(display_freq_10_),
	.datab(display_freq_8_),
	.datac(display_freq_9_),
	.datad(display_freq_11_),
	.cin(gnd),
	.combout(hex6_dup0_2_),
	.cout());
// synopsys translate_off
defparam ix8107z52923.lut_mask = 16'hA210;
defparam ix8107z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y23_N22
cycloneii_lcell_comb ix7110z52923(
// Equation(s):
// hex6_dup0_3_ = display_freq_8_ & (display_freq_10_ $ !display_freq_9_) # !display_freq_8_ & (display_freq_10_ & !display_freq_9_ & !display_freq_11_ # !display_freq_10_ & display_freq_9_ & display_freq_11_)

	.dataa(display_freq_10_),
	.datab(display_freq_8_),
	.datac(display_freq_9_),
	.datad(display_freq_11_),
	.cin(gnd),
	.combout(hex6_dup0_3_),
	.cout());
// synopsys translate_off
defparam ix7110z52923.lut_mask = 16'h9486;
defparam ix7110z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y23_N16
cycloneii_lcell_comb ix6113z52923(
// Equation(s):
// hex6_dup0_4_ = display_freq_9_ & (display_freq_8_ & !display_freq_11_) # !display_freq_9_ & (display_freq_10_ & (!display_freq_11_) # !display_freq_10_ & display_freq_8_)

	.dataa(display_freq_10_),
	.datab(display_freq_8_),
	.datac(display_freq_9_),
	.datad(display_freq_11_),
	.cin(gnd),
	.combout(hex6_dup0_4_),
	.cout());
// synopsys translate_off
defparam ix6113z52923.lut_mask = 16'h04CE;
defparam ix6113z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y23_N26
cycloneii_lcell_comb ix5116z52923(
// Equation(s):
// hex6_dup0_5_ = display_freq_10_ & display_freq_8_ & (display_freq_9_ $ display_freq_11_) # !display_freq_10_ & !display_freq_11_ & (display_freq_8_ # display_freq_9_)

	.dataa(display_freq_10_),
	.datab(display_freq_8_),
	.datac(display_freq_9_),
	.datad(display_freq_11_),
	.cin(gnd),
	.combout(hex6_dup0_5_),
	.cout());
// synopsys translate_off
defparam ix5116z52923.lut_mask = 16'h08D4;
defparam ix5116z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X1_Y23_N12
cycloneii_lcell_comb ix4119z52923(
// Equation(s):
// hex6_dup0_6_ = display_freq_8_ & !display_freq_11_ & (display_freq_10_ $ !display_freq_9_) # !display_freq_8_ & !display_freq_9_ & (display_freq_10_ $ !display_freq_11_)

	.dataa(display_freq_10_),
	.datab(display_freq_8_),
	.datac(display_freq_9_),
	.datad(display_freq_11_),
	.cin(gnd),
	.combout(hex6_dup0_6_),
	.cout());
// synopsys translate_off
defparam ix4119z52923.lut_mask = 16'h0285;
defparam ix4119z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X31_Y14_N28
cycloneii_lcell_comb ix17637z52924(
// Equation(s):
// nx17637z1 = \sw~combout [3] & (\sw~combout [1] # \sw~combout [0] # \sw~combout [2])

	.dataa(\sw~combout [1]),
	.datab(\sw~combout [0]),
	.datac(\sw~combout [3]),
	.datad(\sw~combout [2]),
	.cin(gnd),
	.combout(nx17637z1),
	.cout());
// synopsys translate_off
defparam ix17637z52924.lut_mask = 16'hF0E0;
defparam ix17637z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X28_Y14_N22
cycloneii_lcell_comb ix17637z52923(
// Equation(s):
// hex7_dup0_0_ = \sw~combout [5] & nx4119z4 & (nx17637z1 # \sw~combout [4])

	.dataa(nx17637z1),
	.datab(\sw~combout [5]),
	.datac(\sw~combout [4]),
	.datad(nx4119z4),
	.cin(gnd),
	.combout(hex7_dup0_0_),
	.cout());
// synopsys translate_off
defparam ix17637z52923.lut_mask = 16'hC800;
defparam ix17637z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at PIN_D13
cycloneii_io clock_27_ibuf(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\clock_27~combout ),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(clock_27));
// synopsys translate_off
defparam clock_27_ibuf.input_async_reset = "none";
defparam clock_27_ibuf.input_power_up = "low";
defparam clock_27_ibuf.input_register_mode = "none";
defparam clock_27_ibuf.input_sync_reset = "none";
defparam clock_27_ibuf.oe_async_reset = "none";
defparam clock_27_ibuf.oe_power_up = "low";
defparam clock_27_ibuf.oe_register_mode = "none";
defparam clock_27_ibuf.oe_sync_reset = "none";
defparam clock_27_ibuf.operation_mode = "input";
defparam clock_27_ibuf.output_async_reset = "none";
defparam clock_27_ibuf.output_power_up = "low";
defparam clock_27_ibuf.output_register_mode = "none";
defparam clock_27_ibuf.output_sync_reset = "none";
// synopsys translate_on

// atom is at PLL_3
cycloneii_pll \u_audio_dac_p1_altpll|pll (
	.ena(vcc),
	.clkswitch(gnd),
	.areset(gnd),
	.pfdena(vcc),
	.testclearlock(gnd),
	.sbdin(gnd),
	.inclk({gnd,\clock_27~combout }),
	.locked(),
	.testupout(),
	.testdownout(),
	.sbdout(),
	.clk(\u_audio_dac_p1_altpll|pll_CLK_bus ));
// synopsys translate_off
defparam \u_audio_dac_p1_altpll|pll .bandwidth = 0;
defparam \u_audio_dac_p1_altpll|pll .bandwidth_type = "auto";
defparam \u_audio_dac_p1_altpll|pll .c0_high = 15;
defparam \u_audio_dac_p1_altpll|pll .c0_initial = 1;
defparam \u_audio_dac_p1_altpll|pll .c0_low = 15;
defparam \u_audio_dac_p1_altpll|pll .c0_mode = "even";
defparam \u_audio_dac_p1_altpll|pll .c0_ph = 0;
defparam \u_audio_dac_p1_altpll|pll .c1_mode = "bypass";
defparam \u_audio_dac_p1_altpll|pll .c1_ph = 0;
defparam \u_audio_dac_p1_altpll|pll .c2_mode = "bypass";
defparam \u_audio_dac_p1_altpll|pll .c2_ph = 0;
defparam \u_audio_dac_p1_altpll|pll .charge_pump_current = 80;
defparam \u_audio_dac_p1_altpll|pll .clk0_duty_cycle = 50;
defparam \u_audio_dac_p1_altpll|pll .clk0_phase_shift = "0";
defparam \u_audio_dac_p1_altpll|pll .clk1_counter = "c0";
defparam \u_audio_dac_p1_altpll|pll .clk1_divide_by = 3;
defparam \u_audio_dac_p1_altpll|pll .clk1_duty_cycle = 50;
defparam \u_audio_dac_p1_altpll|pll .clk1_multiply_by = 2;
defparam \u_audio_dac_p1_altpll|pll .clk1_phase_shift = "0";
defparam \u_audio_dac_p1_altpll|pll .clk2_duty_cycle = 50;
defparam \u_audio_dac_p1_altpll|pll .clk2_phase_shift = "0";
defparam \u_audio_dac_p1_altpll|pll .compensate_clock = "clk1";
defparam \u_audio_dac_p1_altpll|pll .gate_lock_counter = 0;
defparam \u_audio_dac_p1_altpll|pll .gate_lock_signal = "no";
defparam \u_audio_dac_p1_altpll|pll .inclk0_input_frequency = 37037;
defparam \u_audio_dac_p1_altpll|pll .inclk1_input_frequency = 37037;
defparam \u_audio_dac_p1_altpll|pll .invalid_lock_multiplier = 5;
defparam \u_audio_dac_p1_altpll|pll .loop_filter_c = 3;
defparam \u_audio_dac_p1_altpll|pll .loop_filter_r = " 2.500000";
defparam \u_audio_dac_p1_altpll|pll .m = 20;
defparam \u_audio_dac_p1_altpll|pll .m_initial = 1;
defparam \u_audio_dac_p1_altpll|pll .m_ph = 0;
defparam \u_audio_dac_p1_altpll|pll .n = 1;
defparam \u_audio_dac_p1_altpll|pll .operation_mode = "normal";
defparam \u_audio_dac_p1_altpll|pll .pfd_max = 100000;
defparam \u_audio_dac_p1_altpll|pll .pfd_min = 2484;
defparam \u_audio_dac_p1_altpll|pll .pll_compensation_delay = 5840;
defparam \u_audio_dac_p1_altpll|pll .self_reset_on_gated_loss_lock = "off";
defparam \u_audio_dac_p1_altpll|pll .sim_gate_lock_device_behavior = "off";
defparam \u_audio_dac_p1_altpll|pll .simulation_type = "timing";
defparam \u_audio_dac_p1_altpll|pll .valid_lock_multiplier = 1;
defparam \u_audio_dac_p1_altpll|pll .vco_center = 1333;
defparam \u_audio_dac_p1_altpll|pll .vco_max = 2000;
defparam \u_audio_dac_p1_altpll|pll .vco_min = 1000;
// synopsys translate_on

// atom is at CLKCTRL_G11
cycloneii_clkctrl \u_audio_dac_p1_altpll|_clk1~clkctrl (
	.ena(vcc),
	.inclk({gnd,gnd,gnd,\u_audio_dac_p1_altpll|_clk1 }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ));
// synopsys translate_off
defparam \u_audio_dac_p1_altpll|_clk1~clkctrl .clock_type = "global clock";
defparam \u_audio_dac_p1_altpll|_clk1~clkctrl .ena_register_mode = "falling edge";
// synopsys translate_on

// atom is at LCCOMB_X34_Y14_N12
cycloneii_lcell_comb ix51811z52923(
// Equation(s):
// NOT_bit_position_0_ = !bit_position_0_

	.dataa(vcc),
	.datab(vcc),
	.datac(bit_position_0_),
	.datad(vcc),
	.cin(gnd),
	.combout(NOT_bit_position_0_),
	.cout());
// synopsys translate_off
defparam ix51811z52923.lut_mask = 16'h0F0F;
defparam ix51811z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y14_N13
cycloneii_lcell_ff modgen_counter_bit_position_reg_q_0_(
	.clk(\aud_bclk_dup0~clkctrl_outclk ),
	.datain(NOT_bit_position_0_),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(bit_position_0_));

// atom is at LCCOMB_X35_Y14_N22
cycloneii_lcell_comb ix49817z52923(
// Equation(s):
// nx49817z1 = bit_position_2_ $ (bit_position_1_ & bit_position_0_)

	.dataa(bit_position_1_),
	.datab(vcc),
	.datac(bit_position_2_),
	.datad(bit_position_0_),
	.cin(gnd),
	.combout(nx49817z1),
	.cout());
// synopsys translate_off
defparam ix49817z52923.lut_mask = 16'h5AF0;
defparam ix49817z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X35_Y14_N23
cycloneii_lcell_ff modgen_counter_bit_position_reg_q_2_(
	.clk(\aud_bclk_dup0~clkctrl_outclk ),
	.datain(nx49817z1),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(bit_position_2_));

// atom is at LCCOMB_X35_Y14_N16
cycloneii_lcell_comb ix48820z52923(
// Equation(s):
// nx48820z1 = bit_position_3_ $ (bit_position_1_ & bit_position_2_ & bit_position_0_)

	.dataa(bit_position_1_),
	.datab(bit_position_2_),
	.datac(bit_position_3_),
	.datad(bit_position_0_),
	.cin(gnd),
	.combout(nx48820z1),
	.cout());
// synopsys translate_off
defparam ix48820z52923.lut_mask = 16'h78F0;
defparam ix48820z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X35_Y14_N17
cycloneii_lcell_ff modgen_counter_bit_position_reg_q_3_(
	.clk(\aud_bclk_dup0~clkctrl_outclk ),
	.datain(nx48820z1),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(bit_position_3_));

// atom is at LCCOMB_X33_Y2_N14
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52931 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx52268z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z15  & !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z16  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z15  & 
// (\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z16  # GND)
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z14  = CARRY(!\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z16  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z15 )

	.dataa(vcc),
	.datab(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z15 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z16 ),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx52268z1 ),
	.cout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z14 ));
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52931 .lut_mask = 16'h3C3F;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at PIN_G26
cycloneii_io key_ibuf_0_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\key~combout [0]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(key[0]));
// synopsys translate_off
defparam key_ibuf_0_.input_async_reset = "none";
defparam key_ibuf_0_.input_power_up = "low";
defparam key_ibuf_0_.input_register_mode = "none";
defparam key_ibuf_0_.input_sync_reset = "none";
defparam key_ibuf_0_.oe_async_reset = "none";
defparam key_ibuf_0_.oe_power_up = "low";
defparam key_ibuf_0_.oe_register_mode = "none";
defparam key_ibuf_0_.oe_sync_reset = "none";
defparam key_ibuf_0_.operation_mode = "input";
defparam key_ibuf_0_.output_async_reset = "none";
defparam key_ibuf_0_.output_power_up = "low";
defparam key_ibuf_0_.output_register_mode = "none";
defparam key_ibuf_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at LCCOMB_X34_Y2_N30
cycloneii_lcell_comb ix48238z52923(
// Equation(s):
// nx48238z1 = !\key~combout [0] # !nx50205z2

	.dataa(vcc),
	.datab(nx50205z2),
	.datac(vcc),
	.datad(\key~combout [0]),
	.cin(gnd),
	.combout(nx48238z1),
	.cout());
// synopsys translate_off
defparam ix48238z52923.lut_mask = 16'h33FF;
defparam ix48238z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X33_Y2_N15
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_1_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx52268z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z15 ));

// atom is at LCCOMB_X33_Y2_N18
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52929 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx54262z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z11  & !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z12  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z11  & 
// (\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z12  # GND)
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z10  = CARRY(!\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z12  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z11 )

	.dataa(vcc),
	.datab(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z11 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z12 ),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx54262z1 ),
	.cout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z10 ));
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52929 .lut_mask = 16'h3C3F;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X33_Y2_N19
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_3_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx54262z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z11 ));

// atom is at LCCOMB_X33_Y2_N22
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52927 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx56256z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z7  & !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z8  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z7  & 
// (\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z8  # GND)
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z6  = CARRY(!\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z8  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z7 )

	.dataa(vcc),
	.datab(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z7 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z8 ),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx56256z1 ),
	.cout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z6 ));
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52927 .lut_mask = 16'h3C3F;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X33_Y2_N23
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_5_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx56256z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z7 ));

// atom is at LCCOMB_X33_Y2_N24
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52926 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx57253z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z5  & (\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z6  $ GND) # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z5  & 
// !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z6  & VCC
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z4  = CARRY(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z5  & !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z6 )

	.dataa(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z5 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z6 ),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx57253z1 ),
	.cout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z4 ));
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52926 .lut_mask = 16'hA50A;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X33_Y2_N25
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_6_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx57253z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z5 ));

// atom is at LCCOMB_X33_Y2_N26
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52925 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx58250z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z3  & !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z4  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z3  & 
// (\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z4  # GND)
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z2  = CARRY(!\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z4  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z3 )

	.dataa(vcc),
	.datab(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z3 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z4 ),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx58250z1 ),
	.cout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z2 ));
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52925 .lut_mask = 16'h3C3F;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X33_Y2_N27
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_7_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx58250z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z3 ));

// atom is at LCCOMB_X33_Y2_N28
cycloneii_lcell_comb \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52923 (
// Equation(s):
// \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z1  = \u_audio_dac_modgen_counter_lrck_1x_div|nx59247z2  $ !\u_audio_dac_modgen_counter_lrck_1x_div|nx2038z1 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_audio_dac_modgen_counter_lrck_1x_div|nx2038z1 ),
	.cin(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z2 ),
	.combout(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z1 ),
	.cout());
// synopsys translate_off
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52923 .lut_mask = 16'hF00F;
defparam \u_audio_dac_modgen_counter_lrck_1x_div|ix59247z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X33_Y2_N29
cycloneii_lcell_ff \u_audio_dac_modgen_counter_lrck_1x_div|reg_q_8_ (
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(nx48238z1),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_audio_dac_modgen_counter_lrck_1x_div|nx2038z1 ));

// atom is at LCCOMB_X34_Y2_N2
cycloneii_lcell_comb ix50205z52924(
// Equation(s):
// nx50205z2 = !\u_audio_dac_modgen_counter_lrck_1x_div|nx2038z1  & (nx50205z3 & !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z5  # !\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z3 )

	.dataa(nx50205z3),
	.datab(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z5 ),
	.datac(\u_audio_dac_modgen_counter_lrck_1x_div|nx2038z1 ),
	.datad(\u_audio_dac_modgen_counter_lrck_1x_div|nx59247z3 ),
	.cin(gnd),
	.combout(nx50205z2),
	.cout());
// synopsys translate_off
defparam ix50205z52924.lut_mask = 16'h020F;
defparam ix50205z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X34_Y2_N28
cycloneii_lcell_comb ix50205z52923(
// Equation(s):
// nx50205z1 = aud_adclrck_dup0 $ !nx50205z2

	.dataa(vcc),
	.datab(vcc),
	.datac(aud_adclrck_dup0),
	.datad(nx50205z2),
	.cin(gnd),
	.combout(nx50205z1),
	.cout());
// synopsys translate_off
defparam ix50205z52923.lut_mask = 16'hF00F;
defparam ix50205z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y2_N29
cycloneii_lcell_ff u_audio_dac_reg_lrck_1x(
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(nx50205z1),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(!\key~combout [0]),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(aud_adclrck_dup0));

// atom is at CLKCTRL_G12
cycloneii_clkctrl \aud_adclrck_dup0~clkctrl (
	.ena(vcc),
	.inclk({gnd,gnd,gnd,aud_adclrck_dup0}),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\aud_adclrck_dup0~clkctrl_outclk ));
// synopsys translate_off
defparam \aud_adclrck_dup0~clkctrl .clock_type = "global clock";
defparam \aud_adclrck_dup0~clkctrl .ena_register_mode = "falling edge";
// synopsys translate_on

// atom is at LCFF_X27_Y14_N13
cycloneii_lcell_ff u_sine_reg_address_3_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx40964z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_3_));

// atom is at LCCOMB_X27_Y14_N8
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52931 (
// Equation(s):
// \u_sine_address_add9_0i1|nx38970z1  = \sw~combout [1] & (u_sine_address_1_ & \u_sine_address_add9_0i1|nx45949z23  & VCC # !u_sine_address_1_ & !\u_sine_address_add9_0i1|nx45949z23 ) # !\sw~combout [1] & (u_sine_address_1_ & 
// !\u_sine_address_add9_0i1|nx45949z23  # !u_sine_address_1_ & (\u_sine_address_add9_0i1|nx45949z23  # GND))
// \u_sine_address_add9_0i1|nx45949z20  = CARRY(\sw~combout [1] & !u_sine_address_1_ & !\u_sine_address_add9_0i1|nx45949z23  # !\sw~combout [1] & (!\u_sine_address_add9_0i1|nx45949z23  # !u_sine_address_1_))

	.dataa(\sw~combout [1]),
	.datab(u_sine_address_1_),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_sine_address_add9_0i1|nx45949z23 ),
	.combout(\u_sine_address_add9_0i1|nx38970z1 ),
	.cout(\u_sine_address_add9_0i1|nx45949z20 ));
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52931 .lut_mask = 16'h9617;
defparam \u_sine_address_add9_0i1|ix45949z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y14_N9
cycloneii_lcell_ff u_sine_reg_address_1_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx38970z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_1_));

// atom is at LCCOMB_X27_Y14_N10
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52930 (
// Equation(s):
// \u_sine_address_add9_0i1|nx39967z1  = (\sw~combout [2] $ u_sine_address_2_ $ !\u_sine_address_add9_0i1|nx45949z20 ) # GND
// \u_sine_address_add9_0i1|nx45949z17  = CARRY(\sw~combout [2] & (u_sine_address_2_ # !\u_sine_address_add9_0i1|nx45949z20 ) # !\sw~combout [2] & u_sine_address_2_ & !\u_sine_address_add9_0i1|nx45949z20 )

	.dataa(\sw~combout [2]),
	.datab(u_sine_address_2_),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_sine_address_add9_0i1|nx45949z20 ),
	.combout(\u_sine_address_add9_0i1|nx39967z1 ),
	.cout(\u_sine_address_add9_0i1|nx45949z17 ));
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52930 .lut_mask = 16'h698E;
defparam \u_sine_address_add9_0i1|ix45949z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y14_N11
cycloneii_lcell_ff u_sine_reg_address_2_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx39967z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_2_));

// atom is at LCCOMB_X27_Y14_N12
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52929 (
// Equation(s):
// \u_sine_address_add9_0i1|nx40964z1  = \sw~combout [3] & (u_sine_address_3_ & \u_sine_address_add9_0i1|nx45949z17  & VCC # !u_sine_address_3_ & !\u_sine_address_add9_0i1|nx45949z17 ) # !\sw~combout [3] & (u_sine_address_3_ & 
// !\u_sine_address_add9_0i1|nx45949z17  # !u_sine_address_3_ & (\u_sine_address_add9_0i1|nx45949z17  # GND))
// \u_sine_address_add9_0i1|nx45949z14  = CARRY(\sw~combout [3] & !u_sine_address_3_ & !\u_sine_address_add9_0i1|nx45949z17  # !\sw~combout [3] & (!\u_sine_address_add9_0i1|nx45949z17  # !u_sine_address_3_))

	.dataa(\sw~combout [3]),
	.datab(u_sine_address_3_),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_sine_address_add9_0i1|nx45949z17 ),
	.combout(\u_sine_address_add9_0i1|nx40964z1 ),
	.cout(\u_sine_address_add9_0i1|nx45949z14 ));
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52929 .lut_mask = 16'h9617;
defparam \u_sine_address_add9_0i1|ix45949z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N14
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52928 (
// Equation(s):
// \u_sine_address_add9_0i1|nx41961z1  = (u_sine_address_4_ $ \sw~combout [4] $ !\u_sine_address_add9_0i1|nx45949z14 ) # GND
// \u_sine_address_add9_0i1|nx45949z11  = CARRY(u_sine_address_4_ & (\sw~combout [4] # !\u_sine_address_add9_0i1|nx45949z14 ) # !u_sine_address_4_ & \sw~combout [4] & !\u_sine_address_add9_0i1|nx45949z14 )

	.dataa(u_sine_address_4_),
	.datab(\sw~combout [4]),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_sine_address_add9_0i1|nx45949z14 ),
	.combout(\u_sine_address_add9_0i1|nx41961z1 ),
	.cout(\u_sine_address_add9_0i1|nx45949z11 ));
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52928 .lut_mask = 16'h698E;
defparam \u_sine_address_add9_0i1|ix45949z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N16
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52927 (
// Equation(s):
// \u_sine_address_add9_0i1|nx42958z1  = u_sine_address_5_ & (\sw~combout [5] & \u_sine_address_add9_0i1|nx45949z11  & VCC # !\sw~combout [5] & !\u_sine_address_add9_0i1|nx45949z11 ) # !u_sine_address_5_ & (\sw~combout [5] & 
// !\u_sine_address_add9_0i1|nx45949z11  # !\sw~combout [5] & (\u_sine_address_add9_0i1|nx45949z11  # GND))
// \u_sine_address_add9_0i1|nx45949z8  = CARRY(u_sine_address_5_ & !\sw~combout [5] & !\u_sine_address_add9_0i1|nx45949z11  # !u_sine_address_5_ & (!\u_sine_address_add9_0i1|nx45949z11  # !\sw~combout [5]))

	.dataa(u_sine_address_5_),
	.datab(\sw~combout [5]),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_sine_address_add9_0i1|nx45949z11 ),
	.combout(\u_sine_address_add9_0i1|nx42958z1 ),
	.cout(\u_sine_address_add9_0i1|nx45949z8 ));
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52927 .lut_mask = 16'h9617;
defparam \u_sine_address_add9_0i1|ix45949z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y14_N19
cycloneii_lcell_ff u_sine_reg_address_6_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx43955z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_6_));

// atom is at LCCOMB_X27_Y14_N18
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52926 (
// Equation(s):
// \u_sine_address_add9_0i1|nx43955z1  = (\sw~combout [6] $ u_sine_address_6_ $ !\u_sine_address_add9_0i1|nx45949z8 ) # GND
// \u_sine_address_add9_0i1|nx45949z5  = CARRY(\sw~combout [6] & (u_sine_address_6_ # !\u_sine_address_add9_0i1|nx45949z8 ) # !\sw~combout [6] & u_sine_address_6_ & !\u_sine_address_add9_0i1|nx45949z8 )

	.dataa(\sw~combout [6]),
	.datab(u_sine_address_6_),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_sine_address_add9_0i1|nx45949z8 ),
	.combout(\u_sine_address_add9_0i1|nx43955z1 ),
	.cout(\u_sine_address_add9_0i1|nx45949z5 ));
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52926 .lut_mask = 16'h698E;
defparam \u_sine_address_add9_0i1|ix45949z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X27_Y14_N20
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52925 (
// Equation(s):
// \u_sine_address_add9_0i1|nx44952z1  = u_sine_address_7_ & !\u_sine_address_add9_0i1|nx45949z5  # !u_sine_address_7_ & (\u_sine_address_add9_0i1|nx45949z5  # GND)
// \u_sine_address_add9_0i1|nx45949z3  = CARRY(!\u_sine_address_add9_0i1|nx45949z5  # !u_sine_address_7_)

	.dataa(u_sine_address_7_),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_sine_address_add9_0i1|nx45949z5 ),
	.combout(\u_sine_address_add9_0i1|nx44952z1 ),
	.cout(\u_sine_address_add9_0i1|nx45949z3 ));
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52925 .lut_mask = 16'h5A5F;
defparam \u_sine_address_add9_0i1|ix45949z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y14_N23
cycloneii_lcell_ff u_sine_reg_address_8_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_sine_address_add9_0i1|nx45949z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_sine_address_8_));

// atom is at LCCOMB_X27_Y14_N22
cycloneii_lcell_comb \u_sine_address_add9_0i1|ix45949z52923 (
// Equation(s):
// \u_sine_address_add9_0i1|nx45949z1  = \u_sine_address_add9_0i1|nx45949z3  $ !u_sine_address_8_

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(u_sine_address_8_),
	.cin(\u_sine_address_add9_0i1|nx45949z3 ),
	.combout(\u_sine_address_add9_0i1|nx45949z1 ),
	.cout());
// synopsys translate_off
defparam \u_sine_address_add9_0i1|ix45949z52923 .lut_mask = 16'hF00F;
defparam \u_sine_address_add9_0i1|ix45949z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X27_Y16_N6
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52933 (
// Equation(s):
// \u_noise_modgen_counter_address|nx51271z1  = \u_noise_modgen_counter_address|q_0_  $ VCC
// \u_noise_modgen_counter_address|nx60244z10  = CARRY(\u_noise_modgen_counter_address|q_0_ )

	.dataa(\u_noise_modgen_counter_address|q_0_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_noise_modgen_counter_address|nx51271z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z10 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52933 .lut_mask = 16'h55AA;
defparam \u_noise_modgen_counter_address|ix60244z52933 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N7
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx51271z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_0_ ));

// atom is at LCCOMB_X27_Y16_N8
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52932 (
// Equation(s):
// \u_noise_modgen_counter_address|nx52268z1  = \u_noise_modgen_counter_address|q_1_  & !\u_noise_modgen_counter_address|nx60244z10  # !\u_noise_modgen_counter_address|q_1_  & (\u_noise_modgen_counter_address|nx60244z10  # GND)
// \u_noise_modgen_counter_address|nx60244z9  = CARRY(!\u_noise_modgen_counter_address|nx60244z10  # !\u_noise_modgen_counter_address|q_1_ )

	.dataa(vcc),
	.datab(\u_noise_modgen_counter_address|q_1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z10 ),
	.combout(\u_noise_modgen_counter_address|nx52268z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z9 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52932 .lut_mask = 16'h3C3F;
defparam \u_noise_modgen_counter_address|ix60244z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N9
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx52268z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_1_ ));

// atom is at LCCOMB_X27_Y16_N10
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52931 (
// Equation(s):
// \u_noise_modgen_counter_address|nx53265z1  = \u_noise_modgen_counter_address|q_2_  & (\u_noise_modgen_counter_address|nx60244z9  $ GND) # !\u_noise_modgen_counter_address|q_2_  & !\u_noise_modgen_counter_address|nx60244z9  & VCC
// \u_noise_modgen_counter_address|nx60244z8  = CARRY(\u_noise_modgen_counter_address|q_2_  & !\u_noise_modgen_counter_address|nx60244z9 )

	.dataa(\u_noise_modgen_counter_address|q_2_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z9 ),
	.combout(\u_noise_modgen_counter_address|nx53265z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z8 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52931 .lut_mask = 16'hA50A;
defparam \u_noise_modgen_counter_address|ix60244z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N11
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx53265z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_2_ ));

// atom is at LCCOMB_X27_Y16_N12
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52930 (
// Equation(s):
// \u_noise_modgen_counter_address|nx54262z1  = \u_noise_modgen_counter_address|q_3_  & !\u_noise_modgen_counter_address|nx60244z8  # !\u_noise_modgen_counter_address|q_3_  & (\u_noise_modgen_counter_address|nx60244z8  # GND)
// \u_noise_modgen_counter_address|nx60244z7  = CARRY(!\u_noise_modgen_counter_address|nx60244z8  # !\u_noise_modgen_counter_address|q_3_ )

	.dataa(\u_noise_modgen_counter_address|q_3_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z8 ),
	.combout(\u_noise_modgen_counter_address|nx54262z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z7 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52930 .lut_mask = 16'h5A5F;
defparam \u_noise_modgen_counter_address|ix60244z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N13
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx54262z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_3_ ));

// atom is at LCCOMB_X27_Y16_N14
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52929 (
// Equation(s):
// \u_noise_modgen_counter_address|nx55259z1  = \u_noise_modgen_counter_address|q_4_  & (\u_noise_modgen_counter_address|nx60244z7  $ GND) # !\u_noise_modgen_counter_address|q_4_  & !\u_noise_modgen_counter_address|nx60244z7  & VCC
// \u_noise_modgen_counter_address|nx60244z6  = CARRY(\u_noise_modgen_counter_address|q_4_  & !\u_noise_modgen_counter_address|nx60244z7 )

	.dataa(vcc),
	.datab(\u_noise_modgen_counter_address|q_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z7 ),
	.combout(\u_noise_modgen_counter_address|nx55259z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z6 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52929 .lut_mask = 16'hC30C;
defparam \u_noise_modgen_counter_address|ix60244z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N15
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx55259z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_4_ ));

// atom is at LCCOMB_X27_Y16_N16
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52928 (
// Equation(s):
// \u_noise_modgen_counter_address|nx56256z1  = \u_noise_modgen_counter_address|q_5_  & !\u_noise_modgen_counter_address|nx60244z6  # !\u_noise_modgen_counter_address|q_5_  & (\u_noise_modgen_counter_address|nx60244z6  # GND)
// \u_noise_modgen_counter_address|nx60244z5  = CARRY(!\u_noise_modgen_counter_address|nx60244z6  # !\u_noise_modgen_counter_address|q_5_ )

	.dataa(\u_noise_modgen_counter_address|q_5_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z6 ),
	.combout(\u_noise_modgen_counter_address|nx56256z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z5 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52928 .lut_mask = 16'h5A5F;
defparam \u_noise_modgen_counter_address|ix60244z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N17
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx56256z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_5_ ));

// atom is at LCCOMB_X27_Y16_N18
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52927 (
// Equation(s):
// \u_noise_modgen_counter_address|nx57253z1  = \u_noise_modgen_counter_address|q_6_  & (\u_noise_modgen_counter_address|nx60244z5  $ GND) # !\u_noise_modgen_counter_address|q_6_  & !\u_noise_modgen_counter_address|nx60244z5  & VCC
// \u_noise_modgen_counter_address|nx60244z4  = CARRY(\u_noise_modgen_counter_address|q_6_  & !\u_noise_modgen_counter_address|nx60244z5 )

	.dataa(vcc),
	.datab(\u_noise_modgen_counter_address|q_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z5 ),
	.combout(\u_noise_modgen_counter_address|nx57253z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z4 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52927 .lut_mask = 16'hC30C;
defparam \u_noise_modgen_counter_address|ix60244z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N19
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx57253z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_6_ ));

// atom is at LCCOMB_X27_Y16_N20
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52926 (
// Equation(s):
// \u_noise_modgen_counter_address|nx58250z1  = \u_noise_modgen_counter_address|q_7_  & !\u_noise_modgen_counter_address|nx60244z4  # !\u_noise_modgen_counter_address|q_7_  & (\u_noise_modgen_counter_address|nx60244z4  # GND)
// \u_noise_modgen_counter_address|nx60244z3  = CARRY(!\u_noise_modgen_counter_address|nx60244z4  # !\u_noise_modgen_counter_address|q_7_ )

	.dataa(\u_noise_modgen_counter_address|q_7_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z4 ),
	.combout(\u_noise_modgen_counter_address|nx58250z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z3 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52926 .lut_mask = 16'h5A5F;
defparam \u_noise_modgen_counter_address|ix60244z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N21
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx58250z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_7_ ));

// atom is at LCCOMB_X27_Y16_N22
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52925 (
// Equation(s):
// \u_noise_modgen_counter_address|nx59247z1  = \u_noise_modgen_counter_address|q_8_  & (\u_noise_modgen_counter_address|nx60244z3  $ GND) # !\u_noise_modgen_counter_address|q_8_  & !\u_noise_modgen_counter_address|nx60244z3  & VCC
// \u_noise_modgen_counter_address|nx60244z2  = CARRY(\u_noise_modgen_counter_address|q_8_  & !\u_noise_modgen_counter_address|nx60244z3 )

	.dataa(vcc),
	.datab(\u_noise_modgen_counter_address|q_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z3 ),
	.combout(\u_noise_modgen_counter_address|nx59247z1 ),
	.cout(\u_noise_modgen_counter_address|nx60244z2 ));
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52925 .lut_mask = 16'hC30C;
defparam \u_noise_modgen_counter_address|ix60244z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N23
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx59247z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_8_ ));

// atom is at LCCOMB_X27_Y16_N24
cycloneii_lcell_comb \u_noise_modgen_counter_address|ix60244z52923 (
// Equation(s):
// \u_noise_modgen_counter_address|nx60244z1  = \u_noise_modgen_counter_address|q_9_  $ \u_noise_modgen_counter_address|nx60244z2 

	.dataa(\u_noise_modgen_counter_address|q_9_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_noise_modgen_counter_address|nx60244z2 ),
	.combout(\u_noise_modgen_counter_address|nx60244z1 ),
	.cout());
// synopsys translate_off
defparam \u_noise_modgen_counter_address|ix60244z52923 .lut_mask = 16'h5A5A;
defparam \u_noise_modgen_counter_address|ix60244z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X27_Y16_N25
cycloneii_lcell_ff \u_noise_modgen_counter_address|reg_q_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_noise_modgen_counter_address|nx60244z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_noise_modgen_counter_address|q_9_ ));

// atom is at M4K_X26_Y15
cycloneii_ram_block \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 (
	.portawe(gnd),
	.portaaddrstall(gnd),
	.portbrewe(vcc),
	.portbaddrstall(gnd),
	.clk0(\aud_adclrck_dup0~clkctrl_outclk ),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(4'b0000),
	.portaaddr({\u_noise_modgen_counter_address|q_9_ ,\u_noise_modgen_counter_address|q_8_ ,\u_noise_modgen_counter_address|q_7_ ,\u_noise_modgen_counter_address|q_6_ ,\u_noise_modgen_counter_address|q_5_ ,\u_noise_modgen_counter_address|q_4_ ,
\u_noise_modgen_counter_address|q_3_ ,\u_noise_modgen_counter_address|q_2_ ,\u_noise_modgen_counter_address|q_1_ ,\u_noise_modgen_counter_address|q_0_ }),
	.portabyteenamasks(1'b1),
	.portbdatain(4'b0000),
	.portbaddr(10'b0000000000),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4_PORTADATAOUT_bus ),
	.portbdataout());
// synopsys translate_off
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .data_interleave_offset_in_bits = 1;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .data_interleave_width_in_bits = 1;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .init_file = "u_noise_modgen_rom_ix24__altsyncram_8_10_1024_2_0.hex";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .init_file_layout = "port_a";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .logical_ram_name = "altsyncram:u_noise_modgen_rom_ix24__ix62120z34212|altsyncram_9nk2:auto_generated|ALTSYNCRAM";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .operation_mode = "rom";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_address_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_address_width = 10;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_byte_enable_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_byte_enable_clock = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_data_in_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_data_out_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_data_out_clock = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_data_width = 4;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_first_address = 0;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_first_bit_number = 4;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_last_address = 1023;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_logical_ram_depth = 1024;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_logical_ram_width = 8;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_write_enable_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_a_write_enable_clock = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_b_address_width = 10;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .port_b_data_width = 4;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .ram_block_type = "M4K";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .safe_write = "err_on_2clk";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .mem_init1 = 2048'h6441071CC8DE5D70761D40307C107E752202FA68CEC0B138C8C693A73757EDF69A8A86C176B00B9787DCC0627C1F65A7319C05622E092119B1D5452D8906942F7F92155731A79E4E36F3F5B6AB61A527BBB5C112CD5F072CD4462D220F3618913DAC993A0242AB7B5D496579A515B87F2DD7786AEC61308B4035E909993CE60AA55580806C67938C40FE2034BDA36E9E9ED1AC81607B3DD8BD24FBBFCFE232BCE1B3C0B68A82FC38FAE6AF35704AFF0B6A1D875A883C0A3E4A0EFFA5619C9A55D281C6E0DDA905EDBF32F21323736EA9B67BCA0D1AC0194E7E753AB70806122991D4589C802A95807AB8A0FE624BE21DF1638F8C73F865138865965874A357E2;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a4 .mem_init0 = 2048'h005AE5EF060ACA6F8EB5B89C615C6D492EB7690F6CDD613F016E49843E3F6ED75825624789A85C62C6E2B42DEDC438A5BDEEA158314108DC266D0D9C451EE4A14BE43DD77A1879D597ACA2380A0C2230C2B9C9CFCA5DDC9B7104377DE21BED9711BA4C1EE5C9E89FEB990A0B74439663CAB11A1754C3BA781F2D92A83679F7637C35FD108C9FD80F061AED3E7010535EBA9727A7C6DD2223A96A63FB8825464BC6A8356B49090009D2D4D201A983D46801E32A314E2C21C84DC875D7DA7158F9BF816213CFFBAEEDB425DA093514C783D366B31FC4EA19E993B70B47932A50B2459CB6FAA2F809FF22B24DAE9F1DD6F2A6FBFA0D3A4912743C2528C459AC1311;
// synopsys translate_on

// atom is at LCCOMB_X34_Y14_N28
cycloneii_lcell_comb ix45891z52925(
// Equation(s):
// raw_audio_9_ = \sw~combout [17] & (\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [5]) # !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [9]

	.dataa(\sw~combout [17]),
	.datab(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [9]),
	.datac(vcc),
	.datad(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [5]),
	.cin(gnd),
	.combout(raw_audio_9_),
	.cout());
// synopsys translate_off
defparam ix45891z52925.lut_mask = 16'hEE44;
defparam ix45891z52925.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X35_Y14_N14
cycloneii_lcell_comb ix45891z52923(
// Equation(s):
// raw_audio_11_ = \sw~combout [17] & (\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [7]) # !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [11]

	.dataa(\sw~combout [17]),
	.datab(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [11]),
	.datac(vcc),
	.datad(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [7]),
	.cin(gnd),
	.combout(raw_audio_11_),
	.cout());
// synopsys translate_off
defparam ix45891z52923.lut_mask = 16'hEE44;
defparam ix45891z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N19
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_11_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__15_ ));

// atom is at LCFF_X49_Y16_N21
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__15_ ));

// atom is at LCFF_X53_Y15_N19
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_2__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__15_ ));

// atom is at LCFF_X54_Y12_N17
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__15_ ));

// atom is at LCFF_X55_Y12_N25
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__15_ ));

// atom is at LCFF_X56_Y9_N21
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_5__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__15_ ));

// atom is at LCFF_X58_Y9_N21
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__15_ ));

// atom is at LCFF_X59_Y9_N25
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__15_ ));

// atom is at LCFF_X60_Y11_N25
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__15_ ));

// atom is at LCFF_X57_Y11_N21
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__15_ ));

// atom is at LCFF_X56_Y11_N23
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__15_ ));

// atom is at LCFF_X54_Y11_N21
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__15_ ));

// atom is at LCCOMB_X35_Y14_N20
cycloneii_lcell_comb ix45891z52924(
// Equation(s):
// raw_audio_10_ = \sw~combout [17] & (\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [6]) # !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [10]

	.dataa(\sw~combout [17]),
	.datab(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [10]),
	.datac(vcc),
	.datad(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [6]),
	.cin(gnd),
	.combout(raw_audio_10_),
	.cout());
// synopsys translate_off
defparam ix45891z52924.lut_mask = 16'hEE44;
defparam ix45891z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N21
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_10_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__10_ ));

// atom is at LCFF_X49_Y16_N19
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__10_ ));

// atom is at LCCOMB_X53_Y15_N28
cycloneii_lcell_comb \u_fir|taps_3__10_~feeder (
// Equation(s):
// \u_fir|taps_3__10_~feeder_combout  = \u_fir|taps_2__10_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_2__10_ ),
	.cin(gnd),
	.combout(\u_fir|taps_3__10_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_3__10_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_3__10_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X53_Y15_N29
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_3__10_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__10_ ));

// atom is at LCFF_X54_Y12_N15
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__10_ ));

// atom is at LCFF_X55_Y12_N21
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__10_ ));

// atom is at LCFF_X56_Y9_N19
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_5__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__10_ ));

// atom is at LCFF_X58_Y9_N19
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__10_ ));

// atom is at LCFF_X59_Y9_N23
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__10_ ));

// atom is at LCFF_X60_Y11_N23
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__10_ ));

// atom is at LCFF_X57_Y11_N19
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__10_ ));

// atom is at LCFF_X56_Y11_N21
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__10_ ));

// atom is at LCFF_X54_Y11_N19
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__10_ ));

// atom is at LCCOMB_X34_Y14_N22
cycloneii_lcell_comb ix45891z52926(
// Equation(s):
// raw_audio_8_ = \sw~combout [17] & \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [4] # !\sw~combout [17] & (\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [8])

	.dataa(\sw~combout [17]),
	.datab(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [4]),
	.datac(vcc),
	.datad(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [8]),
	.cin(gnd),
	.combout(raw_audio_8_),
	.cout());
// synopsys translate_off
defparam ix45891z52926.lut_mask = 16'hDD88;
defparam ix45891z52926.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N17
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_8_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__8_ ));

// atom is at LCFF_X49_Y16_N15
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__8_ ));

// atom is at LCCOMB_X53_Y16_N10
cycloneii_lcell_comb \u_fir|taps_3__8_~feeder (
// Equation(s):
// \u_fir|taps_3__8_~feeder_combout  = \u_fir|taps_2__8_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_2__8_ ),
	.cin(gnd),
	.combout(\u_fir|taps_3__8_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_3__8_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_3__8_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X53_Y16_N11
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_3__8_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__8_ ));

// atom is at LCFF_X54_Y12_N11
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__8_ ));

// atom is at LCFF_X55_Y12_N17
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__8_ ));

// atom is at LCFF_X56_Y9_N15
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_5__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__8_ ));

// atom is at LCFF_X58_Y9_N15
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__8_ ));

// atom is at LCFF_X59_Y9_N19
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__8_ ));

// atom is at LCFF_X60_Y11_N19
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__8_ ));

// atom is at LCFF_X57_Y11_N15
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__8_ ));

// atom is at LCFF_X56_Y11_N17
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__8_ ));

// atom is at LCFF_X54_Y11_N15
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__8_ ));

// atom is at M4K_X26_Y16
cycloneii_ram_block \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 (
	.portawe(gnd),
	.portaaddrstall(gnd),
	.portbrewe(vcc),
	.portbaddrstall(gnd),
	.clk0(\aud_adclrck_dup0~clkctrl_outclk ),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(4'b0000),
	.portaaddr({\u_noise_modgen_counter_address|q_9_ ,\u_noise_modgen_counter_address|q_8_ ,\u_noise_modgen_counter_address|q_7_ ,\u_noise_modgen_counter_address|q_6_ ,\u_noise_modgen_counter_address|q_5_ ,\u_noise_modgen_counter_address|q_4_ ,
\u_noise_modgen_counter_address|q_3_ ,\u_noise_modgen_counter_address|q_2_ ,\u_noise_modgen_counter_address|q_1_ ,\u_noise_modgen_counter_address|q_0_ }),
	.portabyteenamasks(1'b1),
	.portbdatain(4'b0000),
	.portbaddr(10'b0000000000),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0_PORTADATAOUT_bus ),
	.portbdataout());
// synopsys translate_off
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .init_file = "u_noise_modgen_rom_ix24__altsyncram_8_10_1024_2_0.hex";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .init_file_layout = "port_a";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .logical_ram_name = "altsyncram:u_noise_modgen_rom_ix24__ix62120z34212|altsyncram_9nk2:auto_generated|ALTSYNCRAM";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .operation_mode = "rom";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_address_width = 10;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_byte_enable_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_byte_enable_clock = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_data_in_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_data_width = 4;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_last_address = 1023;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 1024;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_logical_ram_width = 8;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_write_enable_clear = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_a_write_enable_clock = "none";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_b_address_width = 10;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .port_b_data_width = 4;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .ram_block_type = "M4K";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .safe_write = "err_on_2clk";
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .mem_init1 = 2048'h1CCEF41A1BE47B8EC04C69D25338F89DDDA04462E827F38DF7D87736B3517F37C3BD4EEDBC309969D6847E3A8D9E0546A6700407E03FE015782194605E54BF10A4F01C8753EB30F760E7C2D24A7EDA6FA4B976DC7F532C2087A84E230F6D5D48D4C1CAAA053DEDF862AEE36B900FC597EC9508728DBB2580FAA9F43FABC5E761295AD818B8612D2FD3F34DA7548C5291536D48CA1E8177D5E75C234648A6DA3CA9E3C16061B05E2CA80E6F469B2EFF2EE04A8257181E62E221EB472AEB49A47B49A61466F543FDB1D62BB60B4B1039E0888665FA817D9179C09FE07C6AE7B3C0FEED2EDA7B5488906381A0965AA97FB8404A5E545D076319B8A259FDCAAA84FC;
defparam \u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|ram_block1a0 .mem_init0 = 2048'hCEB17C5FD83D7C7B444BC9ABCDF44E371EC0BA3773F455A6F03E3250F1DC94A09F7C8DB510F647126FC270098A4B0210E7421635F860E4C07CABE65604A560AD6538DD9E1BFA6628CA10415295D63B13B1E9E22EC1A27E393203E5B0DA4157A7275CCBCBEC41476D599E9C69E6E044F3710F98C4D4E691B32891AA1F76F7F75DEBF5E3FF7A4677932355ECDD8081CC602CBCB9A92763BAFF43ADA446CFF2AB71845993CABA02645D0CB0BF724914112CC94B90AF9E5446AE795051F5CB6BF2B50AA4581EA2EF8B6A1BC774E848C2BEE93DE4DB7640E2C482DFE54DDF6E9B5ADB87A47F137504B2AD332F5F692F00C5B8C4552DBAF9A05C9ADD576576D9B200FE;
// synopsys translate_on

// atom is at LCCOMB_X34_Y14_N18
cycloneii_lcell_comb ix45891z52927(
// Equation(s):
// raw_audio_7_ = \sw~combout [17] & (\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [3]) # !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [7]

	.dataa(\sw~combout [17]),
	.datab(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [7]),
	.datac(vcc),
	.datad(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [3]),
	.cin(gnd),
	.combout(raw_audio_7_),
	.cout());
// synopsys translate_off
defparam ix45891z52927.lut_mask = 16'hEE44;
defparam ix45891z52927.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N15
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_7_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__7_ ));

// atom is at LCFF_X49_Y16_N13
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__7_ ));

// atom is at LCCOMB_X53_Y15_N30
cycloneii_lcell_comb \u_fir|taps_3__7_~feeder (
// Equation(s):
// \u_fir|taps_3__7_~feeder_combout  = \u_fir|taps_2__7_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_2__7_ ),
	.cin(gnd),
	.combout(\u_fir|taps_3__7_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_3__7_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_3__7_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X53_Y15_N31
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_3__7_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__7_ ));

// atom is at LCFF_X54_Y12_N9
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__7_ ));

// atom is at LCFF_X55_Y12_N19
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__7_ ));

// atom is at LCFF_X56_Y9_N13
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_5__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__7_ ));

// atom is at LCFF_X58_Y9_N13
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__7_ ));

// atom is at LCFF_X59_Y9_N17
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__7_ ));

// atom is at LCFF_X60_Y11_N17
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__7_ ));

// atom is at LCFF_X57_Y11_N13
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__7_ ));

// atom is at LCFF_X56_Y11_N15
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__7_ ));

// atom is at LCFF_X54_Y11_N13
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__7_ ));

// atom is at LCCOMB_X34_Y14_N0
cycloneii_lcell_comb ix62120z52923(
// Equation(s):
// raw_audio_5_ = \sw~combout [17] & (\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [1]) # !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [5]

	.dataa(\sw~combout [17]),
	.datab(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [5]),
	.datac(vcc),
	.datad(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [1]),
	.cin(gnd),
	.combout(raw_audio_5_),
	.cout());
// synopsys translate_off
defparam ix62120z52923.lut_mask = 16'hEE44;
defparam ix62120z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N11
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_5_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__5_ ));

// atom is at LCFF_X49_Y16_N9
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__5_ ));

// atom is at LCCOMB_X53_Y16_N0
cycloneii_lcell_comb \u_fir|taps_3__5_~feeder (
// Equation(s):
// \u_fir|taps_3__5_~feeder_combout  = \u_fir|taps_2__5_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_2__5_ ),
	.cin(gnd),
	.combout(\u_fir|taps_3__5_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_3__5_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_3__5_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X53_Y16_N1
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_3__5_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__5_ ));

// atom is at LCFF_X54_Y12_N5
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__5_ ));

// atom is at LCFF_X55_Y12_N15
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__5_ ));

// atom is at LCFF_X56_Y9_N9
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_5__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__5_ ));

// atom is at LCFF_X58_Y9_N9
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__5_ ));

// atom is at LCFF_X59_Y9_N13
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__5_ ));

// atom is at LCFF_X60_Y11_N13
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__5_ ));

// atom is at LCFF_X57_Y11_N9
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__5_ ));

// atom is at LCFF_X56_Y11_N11
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__5_ ));

// atom is at LCFF_X54_Y11_N9
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__5_ ));

// atom is at LCCOMB_X31_Y14_N22
cycloneii_lcell_comb ix45891z52930(
// Equation(s):
// raw_audio_3_ = \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [3] & !\sw~combout [17]

	.dataa(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [3]),
	.datab(\sw~combout [17]),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(raw_audio_3_),
	.cout());
// synopsys translate_off
defparam ix45891z52930.lut_mask = 16'h2222;
defparam ix45891z52930.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N30
cycloneii_lcell_comb \u_fir|taps_1__3_~feeder (
// Equation(s):
// \u_fir|taps_1__3_~feeder_combout  = raw_audio_3_

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(raw_audio_3_),
	.cin(gnd),
	.combout(\u_fir|taps_1__3_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_1__3_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_1__3_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N31
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_1__3_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__3_ ));

// atom is at LCFF_X49_Y16_N5
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__3_ ));

// atom is at LCFF_X53_Y16_N13
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_2__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__3_ ));

// atom is at LCFF_X54_Y12_N1
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__3_ ));

// atom is at LCFF_X55_Y12_N1
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__3_ ));

// atom is at LCCOMB_X56_Y9_N26
cycloneii_lcell_comb \u_fir|taps_6__3_~feeder (
// Equation(s):
// \u_fir|taps_6__3_~feeder_combout  = \u_fir|taps_5__3_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_5__3_ ),
	.cin(gnd),
	.combout(\u_fir|taps_6__3_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_6__3_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_6__3_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X56_Y9_N27
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_6__3_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__3_ ));

// atom is at LCCOMB_X58_Y9_N26
cycloneii_lcell_comb \u_fir|taps_7__3_~feeder (
// Equation(s):
// \u_fir|taps_7__3_~feeder_combout  = \u_fir|taps_6__3_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_6__3_ ),
	.cin(gnd),
	.combout(\u_fir|taps_7__3_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_7__3_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_7__3_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X58_Y9_N27
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_7__3_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__3_ ));

// atom is at LCFF_X59_Y9_N9
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__3_ ));

// atom is at LCFF_X60_Y11_N9
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__3_ ));

// atom is at LCFF_X57_Y11_N5
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__3_ ));

// atom is at LCFF_X56_Y11_N7
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__3_ ));

// atom is at LCFF_X54_Y11_N5
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__3_ ));

// atom is at LCCOMB_X34_Y14_N4
cycloneii_lcell_comb ix45891z52932(
// Equation(s):
// raw_audio_1_ = !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [1]

	.dataa(\sw~combout [17]),
	.datab(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [1]),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(raw_audio_1_),
	.cout());
// synopsys translate_off
defparam ix45891z52932.lut_mask = 16'h4444;
defparam ix45891z52932.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N3
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_1_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__1_ ));

// atom is at LCFF_X49_Y16_N27
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__1_ ));

// atom is at LCFF_X53_Y16_N7
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_2__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__1_ ));

// atom is at LCFF_X53_Y16_N19
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__1_ ));

// atom is at LCCOMB_X55_Y12_N30
cycloneii_lcell_comb \u_fir|taps_5__1_~feeder (
// Equation(s):
// \u_fir|taps_5__1_~feeder_combout  = \u_fir|taps_4__1_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_4__1_ ),
	.cin(gnd),
	.combout(\u_fir|taps_5__1_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_5__1_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_5__1_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X55_Y12_N31
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_5__1_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__1_ ));

// atom is at LCCOMB_X56_Y9_N30
cycloneii_lcell_comb \u_fir|taps_6__1_~feeder (
// Equation(s):
// \u_fir|taps_6__1_~feeder_combout  = \u_fir|taps_5__1_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_5__1_ ),
	.cin(gnd),
	.combout(\u_fir|taps_6__1_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_6__1_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_6__1_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X56_Y9_N31
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_6__1_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__1_ ));

// atom is at LCCOMB_X58_Y9_N30
cycloneii_lcell_comb \u_fir|taps_7__1_~feeder (
// Equation(s):
// \u_fir|taps_7__1_~feeder_combout  = \u_fir|taps_6__1_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_6__1_ ),
	.cin(gnd),
	.combout(\u_fir|taps_7__1_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_7__1_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_7__1_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X58_Y9_N31
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_7__1_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__1_ ));

// atom is at LCFF_X59_Y9_N5
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__1_ ));

// atom is at LCFF_X60_Y11_N5
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__1_ ));

// atom is at LCFF_X57_Y11_N1
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__1_ ));

// atom is at LCFF_X56_Y11_N3
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__1_ ));

// atom is at LCFF_X54_Y11_N1
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__1_ ));

// atom is at LCCOMB_X54_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52940 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z16  = CARRY(\u_fir|taps_12__0_  & \u_fir|taps_12__1_ )

	.dataa(\u_fir|taps_12__0_ ),
	.datab(\u_fir|taps_12__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52940 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52940 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52939 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z15  = CARRY(\u_fir|taps_12__2_  & !\u_fir|taps_12__1_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z16  # !\u_fir|taps_12__2_  & 
// (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z16  # !\u_fir|taps_12__1_ ))

	.dataa(\u_fir|taps_12__2_ ),
	.datab(\u_fir|taps_12__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z16 ),
	.combout(),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z15 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52939 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52939 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52936 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_12__4_  $ \u_fir|taps_12__5_  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z13 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12  = CARRY(\u_fir|taps_12__4_  & (\u_fir|taps_12__5_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z13 ) # !\u_fir|taps_12__4_  & \u_fir|taps_12__5_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z13 )

	.dataa(\u_fir|taps_12__4_ ),
	.datab(\u_fir|taps_12__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z13 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52936 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52935 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_12__6_  & (\u_fir|taps_12__5_  & \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12  & VCC # !\u_fir|taps_12__5_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12 ) # 
// !\u_fir|taps_12__6_  & (\u_fir|taps_12__5_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12  # !\u_fir|taps_12__5_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12  # GND))
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z11  = CARRY(\u_fir|taps_12__6_  & !\u_fir|taps_12__5_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12  # !\u_fir|taps_12__6_  & 
// (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12  # !\u_fir|taps_12__5_ ))

	.dataa(\u_fir|taps_12__6_ ),
	.datab(\u_fir|taps_12__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z12 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52935 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52934 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_12__6_  $ \u_fir|taps_12__7_  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z11 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10  = CARRY(\u_fir|taps_12__6_  & (\u_fir|taps_12__7_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z11 ) # !\u_fir|taps_12__6_  & \u_fir|taps_12__7_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z11 )

	.dataa(\u_fir|taps_12__6_ ),
	.datab(\u_fir|taps_12__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z11 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52934 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52931 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_12__9_  & (\u_fir|taps_12__10_  & \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8  & VCC # !\u_fir|taps_12__10_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8 ) # 
// !\u_fir|taps_12__9_  & (\u_fir|taps_12__10_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8  # !\u_fir|taps_12__10_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8  # GND))
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z7  = CARRY(\u_fir|taps_12__9_  & !\u_fir|taps_12__10_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8  # !\u_fir|taps_12__9_  & 
// (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8  # !\u_fir|taps_12__10_ ))

	.dataa(\u_fir|taps_12__9_ ),
	.datab(\u_fir|taps_12__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z8 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52929 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z6 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|b_10_  = CARRY(\u_fir|taps_12__15_ )

	.dataa(\u_fir|taps_12__15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z6 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|b_10_ ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52929 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_11_ix10225z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|ix10225z52928 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z5  = \u_fir|tap_array_12_filter_block_prod_mults28_0|b_10_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|b_10_ ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z5 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|ix10225z52928 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|ix10225z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X34_Y14_N16
cycloneii_lcell_comb ix45891z52928(
// Equation(s):
// raw_audio_6_ = \sw~combout [17] & (\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [2]) # !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [6]

	.dataa(\sw~combout [17]),
	.datab(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [6]),
	.datac(vcc),
	.datad(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [2]),
	.cin(gnd),
	.combout(raw_audio_6_),
	.cout());
// synopsys translate_off
defparam ix45891z52928.lut_mask = 16'hEE44;
defparam ix45891z52928.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N7
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_6_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__6_ ));

// atom is at LCFF_X49_Y16_N11
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__6_ ));

// atom is at LCCOMB_X53_Y16_N8
cycloneii_lcell_comb \u_fir|taps_3__6_~feeder (
// Equation(s):
// \u_fir|taps_3__6_~feeder_combout  = \u_fir|taps_2__6_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_2__6_ ),
	.cin(gnd),
	.combout(\u_fir|taps_3__6_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_3__6_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_3__6_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X53_Y16_N9
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_3__6_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__6_ ));

// atom is at LCFF_X54_Y12_N7
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__6_ ));

// atom is at LCFF_X55_Y12_N13
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__6_ ));

// atom is at LCFF_X56_Y9_N11
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_5__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__6_ ));

// atom is at LCFF_X58_Y9_N11
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__6_ ));

// atom is at LCFF_X59_Y9_N15
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__6_ ));

// atom is at LCFF_X60_Y11_N15
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__6_ ));

// atom is at LCFF_X57_Y11_N11
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__6_ ));

// atom is at LCFF_X56_Y11_N13
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__6_ ));

// atom is at LCFF_X54_Y11_N11
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__6_ ));

// atom is at LCCOMB_X49_Y16_N28
cycloneii_lcell_comb ix45891z52933(
// Equation(s):
// raw_audio_0_ = !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [0]

	.dataa(\sw~combout [17]),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [0]),
	.cin(gnd),
	.combout(raw_audio_0_),
	.cout());
// synopsys translate_off
defparam ix45891z52933.lut_mask = 16'h5500;
defparam ix45891z52933.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X49_Y16_N29
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_0_),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__0_ ));

// atom is at LCCOMB_X49_Y16_N30
cycloneii_lcell_comb \u_fir|taps_2__0_~feeder (
// Equation(s):
// \u_fir|taps_2__0_~feeder_combout  = \u_fir|taps_1__0_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_1__0_ ),
	.cin(gnd),
	.combout(\u_fir|taps_2__0_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_2__0_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_2__0_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X49_Y16_N31
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_2__0_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__0_ ));

// atom is at LCCOMB_X53_Y16_N2
cycloneii_lcell_comb \u_fir|taps_3__0_~feeder (
// Equation(s):
// \u_fir|taps_3__0_~feeder_combout  = \u_fir|taps_2__0_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_2__0_ ),
	.cin(gnd),
	.combout(\u_fir|taps_3__0_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_3__0_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_3__0_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X53_Y16_N3
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_3__0_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__0_ ));

// atom is at LCFF_X53_Y16_N21
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__0_ ));

// atom is at LCFF_X53_Y16_N17
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__0_ ));

// atom is at LCCOMB_X57_Y9_N28
cycloneii_lcell_comb \u_fir|taps_6__0_~feeder (
// Equation(s):
// \u_fir|taps_6__0_~feeder_combout  = \u_fir|taps_5__0_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_5__0_ ),
	.cin(gnd),
	.combout(\u_fir|taps_6__0_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_6__0_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_6__0_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X57_Y9_N29
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_6__0_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__0_ ));

// atom is at LCFF_X56_Y9_N1
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__0_ ));

// atom is at LCFF_X56_Y9_N3
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__0_ ));

// atom is at LCFF_X56_Y9_N5
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__0_ ));

// atom is at LCCOMB_X60_Y11_N0
cycloneii_lcell_comb \u_fir|taps_10__0_~feeder (
// Equation(s):
// \u_fir|taps_10__0_~feeder_combout  = \u_fir|taps_9__0_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_9__0_ ),
	.cin(gnd),
	.combout(\u_fir|taps_10__0_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_10__0_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_10__0_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X60_Y11_N1
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_10__0_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__0_ ));

// atom is at LCCOMB_X60_Y11_N2
cycloneii_lcell_comb \u_fir|taps_11__0_~feeder (
// Equation(s):
// \u_fir|taps_11__0_~feeder_combout  = \u_fir|taps_10__0_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_10__0_ ),
	.cin(gnd),
	.combout(\u_fir|taps_11__0_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_11__0_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_11__0_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X60_Y11_N3
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_11__0_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__0_ ));

// atom is at LCFF_X53_Y11_N5
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__0_ ));

// atom is at LCCOMB_X53_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52950 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z26  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_2_  & \u_fir|taps_12__0_ )

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_2_ ),
	.datab(\u_fir|taps_12__0_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z26 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52950 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52950 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52949 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z25  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_3_  & !\u_fir|taps_12__1_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z26  # 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_3_  & (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z26  # !\u_fir|taps_12__1_ ))

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_3_ ),
	.datab(\u_fir|taps_12__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z26 ),
	.combout(),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52949 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52949 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52948 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24  = CARRY(\u_fir|taps_12__2_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z25 ) # !\u_fir|taps_12__2_  & 
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z25 )

	.dataa(\u_fir|taps_12__2_ ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z25 ),
	.combout(),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52948 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52948 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52947 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_3__dup_193  = \u_fir|taps_12__3_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_  & \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24  & VCC # 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24 ) # !\u_fir|taps_12__3_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_  & 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24  # GND))
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z23  = CARRY(\u_fir|taps_12__3_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24  # !\u_fir|taps_12__3_  & 
// (!\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_ ))

	.dataa(\u_fir|taps_12__3_ ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z24 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_3__dup_193 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z23 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52947 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52947 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52946 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192  = (\u_fir|taps_12__4_  $ \u_fir|tap_array_12_filter_block_prod_mults28_0|d_6_  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z23 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22  = CARRY(\u_fir|taps_12__4_  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z23 ) # !\u_fir|taps_12__4_  & 
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z23 )

	.dataa(\u_fir|taps_12__4_ ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z23 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52946 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52946 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52944 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8_  $ \u_fir|taps_12__6_  $ !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z21 ) # GND
// \u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8_  & (\u_fir|taps_12__6_  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z21 ) # 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8_  & \u_fir|taps_12__6_  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z21 )

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8_ ),
	.datab(\u_fir|taps_12__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z21 ),
	.combout(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_6__dup_190 ),
	.cout(\u_fir|tap_array_12_filter_block_prod_mults28_0|nx10225z20 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52944 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_prod_mults28_0|modgen_add_12_ix10225z52944 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N13
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_9_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__9_ ));

// atom is at LCFF_X49_Y16_N17
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__9_ ));

// atom is at LCCOMB_X53_Y15_N24
cycloneii_lcell_comb \u_fir|taps_3__9_~feeder (
// Equation(s):
// \u_fir|taps_3__9_~feeder_combout  = \u_fir|taps_2__9_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_2__9_ ),
	.cin(gnd),
	.combout(\u_fir|taps_3__9_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_3__9_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_3__9_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X53_Y15_N25
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_3__9_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__9_ ));

// atom is at LCFF_X54_Y12_N13
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__9_ ));

// atom is at LCFF_X55_Y12_N23
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__9_ ));

// atom is at LCFF_X56_Y9_N17
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_5__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__9_ ));

// atom is at LCFF_X58_Y9_N17
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__9_ ));

// atom is at LCFF_X59_Y9_N21
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__9_ ));

// atom is at LCFF_X60_Y11_N21
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__9_ ));

// atom is at LCFF_X57_Y11_N17
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__9_ ));

// atom is at LCFF_X56_Y11_N19
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__9_ ));

// atom is at LCCOMB_X34_Y14_N2
cycloneii_lcell_comb ix45891z52929(
// Equation(s):
// raw_audio_4_ = \sw~combout [17] & (\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [0]) # !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [4]

	.dataa(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [4]),
	.datab(\u_noise_modgen_rom_ix24__ix62120z34212|auto_generated|q_a [0]),
	.datac(vcc),
	.datad(\sw~combout [17]),
	.cin(gnd),
	.combout(raw_audio_4_),
	.cout());
// synopsys translate_off
defparam ix45891z52929.lut_mask = 16'hCCAA;
defparam ix45891z52929.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N9
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_4_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__4_ ));

// atom is at LCFF_X49_Y16_N7
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__4_ ));

// atom is at LCFF_X53_Y16_N5
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_2__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__4_ ));

// atom is at LCFF_X54_Y12_N3
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__4_ ));

// atom is at LCFF_X55_Y12_N9
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_4__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__4_ ));

// atom is at LCFF_X56_Y9_N7
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_5__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__4_ ));

// atom is at LCFF_X58_Y9_N7
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_6__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__4_ ));

// atom is at LCFF_X59_Y9_N11
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__4_ ));

// atom is at LCFF_X60_Y11_N11
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__4_ ));

// atom is at LCFF_X57_Y11_N7
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__4_ ));

// atom is at LCFF_X56_Y11_N9
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__4_ ));

// atom is at LCCOMB_X34_Y14_N10
cycloneii_lcell_comb ix45891z52931(
// Equation(s):
// raw_audio_2_ = !\sw~combout [17] & \u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [2]

	.dataa(\sw~combout [17]),
	.datab(\u_sine_modgen_rom_ix21__ix62120z58996|auto_generated|q_a [2]),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(raw_audio_2_),
	.cout());
// synopsys translate_off
defparam ix45891z52931.lut_mask = 16'h4444;
defparam ix45891z52931.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X48_Y16_N5
cycloneii_lcell_ff \u_fir|tap_array_1_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(raw_audio_2_),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_1__2_ ));

// atom is at LCFF_X49_Y16_N3
cycloneii_lcell_ff \u_fir|tap_array_2_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_1__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_2__2_ ));

// atom is at LCFF_X53_Y16_N15
cycloneii_lcell_ff \u_fir|tap_array_3_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_2__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_3__2_ ));

// atom is at LCFF_X53_Y16_N23
cycloneii_lcell_ff \u_fir|tap_array_4_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_3__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_4__2_ ));

// atom is at LCCOMB_X55_Y12_N2
cycloneii_lcell_comb \u_fir|taps_5__2_~feeder (
// Equation(s):
// \u_fir|taps_5__2_~feeder_combout  = \u_fir|taps_4__2_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_4__2_ ),
	.cin(gnd),
	.combout(\u_fir|taps_5__2_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_5__2_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_5__2_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X55_Y12_N3
cycloneii_lcell_ff \u_fir|tap_array_5_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_5__2_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_5__2_ ));

// atom is at LCCOMB_X56_Y9_N28
cycloneii_lcell_comb \u_fir|taps_6__2_~feeder (
// Equation(s):
// \u_fir|taps_6__2_~feeder_combout  = \u_fir|taps_5__2_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_5__2_ ),
	.cin(gnd),
	.combout(\u_fir|taps_6__2_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_6__2_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_6__2_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X56_Y9_N29
cycloneii_lcell_ff \u_fir|tap_array_6_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_6__2_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_6__2_ ));

// atom is at LCCOMB_X58_Y9_N28
cycloneii_lcell_comb \u_fir|taps_7__2_~feeder (
// Equation(s):
// \u_fir|taps_7__2_~feeder_combout  = \u_fir|taps_6__2_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_6__2_ ),
	.cin(gnd),
	.combout(\u_fir|taps_7__2_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_7__2_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_7__2_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X58_Y9_N29
cycloneii_lcell_ff \u_fir|tap_array_7_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_7__2_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_7__2_ ));

// atom is at LCFF_X59_Y9_N7
cycloneii_lcell_ff \u_fir|tap_array_8_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_7__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_8__2_ ));

// atom is at LCFF_X60_Y11_N7
cycloneii_lcell_ff \u_fir|tap_array_9_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_8__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_9__2_ ));

// atom is at LCFF_X57_Y11_N3
cycloneii_lcell_ff \u_fir|tap_array_10_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_9__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_10__2_ ));

// atom is at LCFF_X56_Y11_N5
cycloneii_lcell_ff \u_fir|tap_array_11_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_10__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_11__2_ ));

// atom is at LCCOMB_X56_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52936 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z13  = CARRY(\u_fir|taps_11__0_  & \u_fir|taps_11__1_ )

	.dataa(\u_fir|taps_11__0_ ),
	.datab(\u_fir|taps_11__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52935 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z12  = CARRY(\u_fir|taps_11__1_  & !\u_fir|taps_11__2_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_11__1_  & 
// (!\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_11__2_ ))

	.dataa(\u_fir|taps_11__1_ ),
	.datab(\u_fir|taps_11__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z13 ),
	.combout(),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52934 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11  = CARRY(\u_fir|taps_11__3_  & (\u_fir|taps_11__2_  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z12 ) # !\u_fir|taps_11__3_  & \u_fir|taps_11__2_  & 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z12 )

	.dataa(\u_fir|taps_11__3_ ),
	.datab(\u_fir|taps_11__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z12 ),
	.combout(),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52933 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_11__3_  & (\u_fir|taps_11__4_  & \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11  & VCC # !\u_fir|taps_11__4_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11 ) # 
// !\u_fir|taps_11__3_  & (\u_fir|taps_11__4_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_11__4_  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11  # GND))
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z10  = CARRY(\u_fir|taps_11__3_  & !\u_fir|taps_11__4_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_11__3_  & 
// (!\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_11__4_ ))

	.dataa(\u_fir|taps_11__3_ ),
	.datab(\u_fir|taps_11__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z11 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52932 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_11__5_  $ \u_fir|taps_11__4_  $ !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z10 ) # GND
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9  = CARRY(\u_fir|taps_11__5_  & (\u_fir|taps_11__4_  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z10 ) # !\u_fir|taps_11__5_  & \u_fir|taps_11__4_  & 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z10 )

	.dataa(\u_fir|taps_11__5_ ),
	.datab(\u_fir|taps_11__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z10 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52931 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_11__6_  & (\u_fir|taps_11__5_  & \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9  & VCC # !\u_fir|taps_11__5_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9 ) # 
// !\u_fir|taps_11__6_  & (\u_fir|taps_11__5_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_11__5_  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9  # GND))
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z8  = CARRY(\u_fir|taps_11__6_  & !\u_fir|taps_11__5_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_11__6_  & (!\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9  
// # !\u_fir|taps_11__5_ ))

	.dataa(\u_fir|taps_11__6_ ),
	.datab(\u_fir|taps_11__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z9 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52930 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_11__6_  $ \u_fir|taps_11__7_  $ !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z8 ) # GND
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7  = CARRY(\u_fir|taps_11__6_  & (\u_fir|taps_11__7_  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z8 ) # !\u_fir|taps_11__6_  & \u_fir|taps_11__7_  & 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z8 )

	.dataa(\u_fir|taps_11__6_ ),
	.datab(\u_fir|taps_11__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z8 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52928 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_11__8_  $ \u_fir|taps_11__9_  $ !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z6 ) # GND
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5  = CARRY(\u_fir|taps_11__8_  & (\u_fir|taps_11__9_  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z6 ) # !\u_fir|taps_11__8_  & \u_fir|taps_11__9_  & 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z6 )

	.dataa(\u_fir|taps_11__8_ ),
	.datab(\u_fir|taps_11__9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z6 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52927 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_11__10_  & (\u_fir|taps_11__9_  & \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5  & VCC # !\u_fir|taps_11__9_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5 ) # 
// !\u_fir|taps_11__10_  & (\u_fir|taps_11__9_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_11__9_  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5  # GND))
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z4  = CARRY(\u_fir|taps_11__10_  & !\u_fir|taps_11__9_  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_11__10_  & (!\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5 
//  # !\u_fir|taps_11__9_ ))

	.dataa(\u_fir|taps_11__10_ ),
	.datab(\u_fir|taps_11__9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z5 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52926 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_11__10_  $ \u_fir|taps_11__15_  $ !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z4 ) # GND
// \u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z3  = CARRY(\u_fir|taps_11__10_  & (\u_fir|taps_11__15_  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z4 ) # !\u_fir|taps_11__10_  & \u_fir|taps_11__15_  & 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z4 )

	.dataa(\u_fir|taps_11__10_ ),
	.datab(\u_fir|taps_11__15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z4 ),
	.combout(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_11_filter_block_prod_mults28_0|nx9228z3 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52926 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_prod_mults28_0|modgen_add_10_ix9228z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52936 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z13  = CARRY(\u_fir|taps_9__0_  & \u_fir|taps_9__1_ )

	.dataa(\u_fir|taps_9__0_ ),
	.datab(\u_fir|taps_9__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52935 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z12  = CARRY(\u_fir|taps_9__2_  & !\u_fir|taps_9__1_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_9__2_  & (!\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z13  # 
// !\u_fir|taps_9__1_ ))

	.dataa(\u_fir|taps_9__2_ ),
	.datab(\u_fir|taps_9__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z13 ),
	.combout(),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52934 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11  = CARRY(\u_fir|taps_9__2_  & (\u_fir|taps_9__3_  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z12 ) # !\u_fir|taps_9__2_  & \u_fir|taps_9__3_  & 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z12 )

	.dataa(\u_fir|taps_9__2_ ),
	.datab(\u_fir|taps_9__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z12 ),
	.combout(),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52932 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_9__4_  $ \u_fir|taps_9__5_  $ !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z10 ) # GND
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9  = CARRY(\u_fir|taps_9__4_  & (\u_fir|taps_9__5_  # !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z10 ) # !\u_fir|taps_9__4_  & \u_fir|taps_9__5_  & 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z10 )

	.dataa(\u_fir|taps_9__4_ ),
	.datab(\u_fir|taps_9__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z10 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52931 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_9__5_  & (\u_fir|taps_9__6_  & \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9  & VCC # !\u_fir|taps_9__6_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9 ) # 
// !\u_fir|taps_9__5_  & (\u_fir|taps_9__6_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_9__6_  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9  # GND))
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z8  = CARRY(\u_fir|taps_9__5_  & !\u_fir|taps_9__6_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_9__5_  & (!\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9  # 
// !\u_fir|taps_9__6_ ))

	.dataa(\u_fir|taps_9__5_ ),
	.datab(\u_fir|taps_9__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z9 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52929 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_9__7_  & (\u_fir|taps_9__8_  & \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7  & VCC # !\u_fir|taps_9__8_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7 ) # 
// !\u_fir|taps_9__7_  & (\u_fir|taps_9__8_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_9__8_  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7  # GND))
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z6  = CARRY(\u_fir|taps_9__7_  & !\u_fir|taps_9__8_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_9__7_  & (!\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7  # 
// !\u_fir|taps_9__8_ ))

	.dataa(\u_fir|taps_9__7_ ),
	.datab(\u_fir|taps_9__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z7 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N0
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52936 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z13  = CARRY(\u_fir|taps_7__0_  & \u_fir|taps_7__1_ )

	.dataa(\u_fir|taps_7__0_ ),
	.datab(\u_fir|taps_7__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N2
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52935 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z12  = CARRY(\u_fir|taps_7__2_  & !\u_fir|taps_7__1_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_7__2_  & (!\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z13  # 
// !\u_fir|taps_7__1_ ))

	.dataa(\u_fir|taps_7__2_ ),
	.datab(\u_fir|taps_7__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z13 ),
	.combout(),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N4
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52934 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11  = CARRY(\u_fir|taps_7__2_  & (\u_fir|taps_7__3_  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z12 ) # !\u_fir|taps_7__2_  & \u_fir|taps_7__3_  & 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z12 )

	.dataa(\u_fir|taps_7__2_ ),
	.datab(\u_fir|taps_7__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z12 ),
	.combout(),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N6
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52933 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_7__4_  & (\u_fir|taps_7__3_  & \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11  & VCC # !\u_fir|taps_7__3_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11 ) # 
// !\u_fir|taps_7__4_  & (\u_fir|taps_7__3_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_7__3_  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11  # GND))
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z10  = CARRY(\u_fir|taps_7__4_  & !\u_fir|taps_7__3_  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_7__4_  & (!\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11  # 
// !\u_fir|taps_7__3_ ))

	.dataa(\u_fir|taps_7__4_ ),
	.datab(\u_fir|taps_7__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z11 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N8
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52932 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_7__4_  $ \u_fir|taps_7__5_  $ !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z10 ) # GND
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9  = CARRY(\u_fir|taps_7__4_  & (\u_fir|taps_7__5_  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z10 ) # !\u_fir|taps_7__4_  & \u_fir|taps_7__5_  & 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z10 )

	.dataa(\u_fir|taps_7__4_ ),
	.datab(\u_fir|taps_7__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z10 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y9_N12
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52930 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_7__6_  $ \u_fir|taps_7__7_  $ !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z8 ) # GND
// \u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7  = CARRY(\u_fir|taps_7__6_  & (\u_fir|taps_7__7_  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z8 ) # !\u_fir|taps_7__6_  & \u_fir|taps_7__7_  & 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z8 )

	.dataa(\u_fir|taps_7__6_ ),
	.datab(\u_fir|taps_7__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z8 ),
	.combout(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_7_filter_block_prod_mults28_0|nx9228z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_prod_mults28_0|modgen_add_6_ix9228z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N0
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52940 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z16  = CARRY(\u_fir|taps_6__0_  & \u_fir|taps_6__1_ )

	.dataa(\u_fir|taps_6__0_ ),
	.datab(\u_fir|taps_6__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52940 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52940 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N2
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52939 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z15  = CARRY(\u_fir|taps_6__2_  & !\u_fir|taps_6__1_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z16  # !\u_fir|taps_6__2_  & (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z16  
// # !\u_fir|taps_6__1_ ))

	.dataa(\u_fir|taps_6__2_ ),
	.datab(\u_fir|taps_6__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z16 ),
	.combout(),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z15 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52939 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52939 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N6
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52937 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_6__4_  & (\u_fir|taps_6__3_  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14  & VCC # !\u_fir|taps_6__3_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14 ) # 
// !\u_fir|taps_6__4_  & (\u_fir|taps_6__3_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14  # !\u_fir|taps_6__3_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14  # GND))
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z13  = CARRY(\u_fir|taps_6__4_  & !\u_fir|taps_6__3_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14  # !\u_fir|taps_6__4_  & (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14  
// # !\u_fir|taps_6__3_ ))

	.dataa(\u_fir|taps_6__4_ ),
	.datab(\u_fir|taps_6__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z14 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52937 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N14
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52933 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_6__7_  & (\u_fir|taps_6__8_  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10  & VCC # !\u_fir|taps_6__8_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10 ) # 
// !\u_fir|taps_6__7_  & (\u_fir|taps_6__8_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10  # !\u_fir|taps_6__8_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10  # GND))
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z9  = CARRY(\u_fir|taps_6__7_  & !\u_fir|taps_6__8_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10  # !\u_fir|taps_6__7_  & (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10  # 
// !\u_fir|taps_6__8_ ))

	.dataa(\u_fir|taps_6__7_ ),
	.datab(\u_fir|taps_6__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z10 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N0
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52950 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z26  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_2_  & \u_fir|taps_6__0_ )

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_2_ ),
	.datab(\u_fir|taps_6__0_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z26 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52950 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52950 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N2
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52949 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z25  = CARRY(\u_fir|taps_6__1_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_3_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z26  # !\u_fir|taps_6__1_  & 
// (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z26  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_3_ ))

	.dataa(\u_fir|taps_6__1_ ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z26 ),
	.combout(),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52949 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52949 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N4
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52948 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4_  & (\u_fir|taps_6__2_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z25 ) # 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4_  & \u_fir|taps_6__2_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z25 )

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_4_ ),
	.datab(\u_fir|taps_6__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z25 ),
	.combout(),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z24 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52948 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52948 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N10
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52945 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_5__dup_191  = \u_fir|taps_6__5_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22  & VCC # 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22 ) # !\u_fir|taps_6__5_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22 
//  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22  # GND))
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z21  = CARRY(\u_fir|taps_6__5_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22  # !\u_fir|taps_6__5_  & 
// (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_ ))

	.dataa(\u_fir|taps_6__5_ ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z22 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_5__dup_191 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z21 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52945 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52945 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N0
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|taps_4__3_  $ VCC) # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|taps_4__3_  & VCC
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|taps_4__3_ )

	.dataa(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|taps_4__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N2
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|taps_4__4_  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46  & VCC # !\u_fir|taps_4__4_  & 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|taps_4__4_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|taps_4__4_  & 
// (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|taps_4__4_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|taps_4__4_ ))

	.dataa(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|taps_4__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N0
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_5_filter_block_prod_mults28_0|d_3_  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx37973z1  $ VCC) # !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_3_  & 
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx37973z1  & VCC
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_3_  & \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx37973z1 )

	.dataa(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_3_ ),
	.datab(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx37973z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N2
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_5_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46  & VCC # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_4_  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1  & 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46  # GND))
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_4_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46  # 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_4_  & (!\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1 ))

	.dataa(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_4_ ),
	.datab(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx38970z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N4
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|tap_array_6_filter_block_prod_mults28_0|d_5__dup_191  $ !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_5__dup_191  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z43 ) 
// # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|tap_array_6_filter_block_prod_mults28_0|d_5__dup_191  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_5__dup_191 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N6
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_  & \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_  & 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx40964z1  & (!\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_ ))

	.dataa(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx40964z1 ),
	.datab(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N4
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52936 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z13  = CARRY(\u_fir|taps_8__0_  & \u_fir|taps_8__1_ )

	.dataa(\u_fir|taps_8__0_ ),
	.datab(\u_fir|taps_8__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N6
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52935 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z12  = CARRY(\u_fir|taps_8__2_  & !\u_fir|taps_8__1_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_8__2_  & (!\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z13  # 
// !\u_fir|taps_8__1_ ))

	.dataa(\u_fir|taps_8__2_ ),
	.datab(\u_fir|taps_8__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z13 ),
	.combout(),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N8
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52934 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11  = CARRY(\u_fir|taps_8__2_  & (\u_fir|taps_8__3_  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z12 ) # !\u_fir|taps_8__2_  & \u_fir|taps_8__3_  & 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z12 )

	.dataa(\u_fir|taps_8__2_ ),
	.datab(\u_fir|taps_8__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z12 ),
	.combout(),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N10
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52933 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_8__4_  & (\u_fir|taps_8__3_  & \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11  & VCC # !\u_fir|taps_8__3_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11 ) # 
// !\u_fir|taps_8__4_  & (\u_fir|taps_8__3_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_8__3_  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11  # GND))
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z10  = CARRY(\u_fir|taps_8__4_  & !\u_fir|taps_8__3_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11  # !\u_fir|taps_8__4_  & (!\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11  # 
// !\u_fir|taps_8__3_ ))

	.dataa(\u_fir|taps_8__4_ ),
	.datab(\u_fir|taps_8__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z11 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N12
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52932 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_8__5_  $ \u_fir|taps_8__4_  $ !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z10 ) # GND
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9  = CARRY(\u_fir|taps_8__5_  & (\u_fir|taps_8__4_  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z10 ) # !\u_fir|taps_8__5_  & \u_fir|taps_8__4_  & 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z10 )

	.dataa(\u_fir|taps_8__5_ ),
	.datab(\u_fir|taps_8__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z10 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N14
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52931 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_8__5_  & (\u_fir|taps_8__6_  & \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9  & VCC # !\u_fir|taps_8__6_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9 ) # 
// !\u_fir|taps_8__5_  & (\u_fir|taps_8__6_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_8__6_  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9  # GND))
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z8  = CARRY(\u_fir|taps_8__5_  & !\u_fir|taps_8__6_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_8__5_  & (!\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9  # 
// !\u_fir|taps_8__6_ ))

	.dataa(\u_fir|taps_8__5_ ),
	.datab(\u_fir|taps_8__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z9 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N0
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_3_  $ VCC) # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx37973z1  & 
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_3_  & VCC
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|tap_array_8_filter_block_prod_mults28_0|d_3_ )

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N6
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_8_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1  & 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_6_  & (!\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1 ))

	.dataa(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_6_ ),
	.datab(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx40964z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_9_filter_block_prod_mults28_0|d_3_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx37973z1  $ VCC) # !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_3_  & 
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx37973z1  & VCC
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_3_  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx37973z1 )

	.dataa(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_3_ ),
	.datab(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx37973z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_9_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1  & 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_6_  & (!\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1 ))

	.dataa(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_6_ ),
	.datab(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx40964z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|tap_array_9_filter_block_prod_mults28_0|d_7_  $ !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|d_7_  # !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|tap_array_9_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52936 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z13  = CARRY(\u_fir|taps_10__0_  & \u_fir|taps_10__1_ )

	.dataa(\u_fir|taps_10__0_ ),
	.datab(\u_fir|taps_10__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52935 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z12  = CARRY(\u_fir|taps_10__1_  & !\u_fir|taps_10__2_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_10__1_  & 
// (!\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_10__2_ ))

	.dataa(\u_fir|taps_10__1_ ),
	.datab(\u_fir|taps_10__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z13 ),
	.combout(),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52934 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11  = CARRY(\u_fir|taps_10__3_  & (\u_fir|taps_10__2_  # !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z12 ) # !\u_fir|taps_10__3_  & \u_fir|taps_10__2_  & 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z12 )

	.dataa(\u_fir|taps_10__3_ ),
	.datab(\u_fir|taps_10__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z12 ),
	.combout(),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52932 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_10__4_  $ \u_fir|taps_10__5_  $ !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z10 ) # GND
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9  = CARRY(\u_fir|taps_10__4_  & (\u_fir|taps_10__5_  # !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z10 ) # !\u_fir|taps_10__4_  & \u_fir|taps_10__5_  & 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z10 )

	.dataa(\u_fir|taps_10__4_ ),
	.datab(\u_fir|taps_10__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z10 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52931 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_10__6_  & (\u_fir|taps_10__5_  & \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9  & VCC # !\u_fir|taps_10__5_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9 ) # 
// !\u_fir|taps_10__6_  & (\u_fir|taps_10__5_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_10__5_  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9  # GND))
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z8  = CARRY(\u_fir|taps_10__6_  & !\u_fir|taps_10__5_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_10__6_  & (!\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9  
// # !\u_fir|taps_10__5_ ))

	.dataa(\u_fir|taps_10__6_ ),
	.datab(\u_fir|taps_10__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z9 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_10_filter_block_prod_mults28_0|d_7_  $ \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx41961z1  $ !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx41961z1  # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_10_filter_block_prod_mults28_0|d_7_  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx41961z1  & !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx41961z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_10_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|tap_array_11_filter_block_prod_mults28_0|d_5_  $ !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_5_  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|tap_array_11_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_7_  $ \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx41961z1  $ !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx41961z1  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_7_  & \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx41961z1  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx41961z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_  & 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx42958z1  & (!\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_ ))

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx42958z1 ),
	.datab(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx43955z1  $ \u_fir|tap_array_11_filter_block_prod_mults28_0|d_9_  $ !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx43955z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_9_  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx43955z1  & \u_fir|tap_array_11_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx43955z1 ),
	.datab(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_10_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_  & 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx44952z1  & (!\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_ ))

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx44952z1 ),
	.datab(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_11_filter_block_prod_mults28_0|d_11_  $ !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_11_filter_block_prod_mults28_0|d_11_  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_11_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_10_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_11_filter_block_prod_mults28_0|d_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_11_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_3__dup_193  $ VCC) # 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|tap_array_12_filter_block_prod_mults28_0|d_3__dup_193  & VCC
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|tap_array_12_filter_block_prod_mults28_0|d_3__dup_193 )

	.dataa(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_3__dup_193 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N2
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52938 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1  = \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx38970z1  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46  & 
// VCC # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46 ) # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx38970z1  & 
// (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46  
// # GND))
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z43  = CARRY(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx38970z1  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192  & 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx38970z1  & (!\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192 
// ))

	.dataa(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx38970z1 ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_4__dup_192 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z46 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx38970z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z43 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52938 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7__dup_189  $ \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx41961z1  $ !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z37 ) # 
// GND
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7__dup_189  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx41961z1  # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z37 ) # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7__dup_189  & \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx41961z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_7__dup_189 ),
	.datab(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx41961z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_12_filter_block_prod_mults28_0|d_8__dup_188  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34  & 
// VCC # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8__dup_188  & 
// (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34  # 
// GND))
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8__dup_188  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8__dup_188  & (!\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1 
// ))

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_8__dup_188 ),
	.datab(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_12_filter_block_prod_mults28_0|d_10__dup_186  & (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28  & 
// VCC # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10__dup_186  & 
// (\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28  # 
// GND))
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10__dup_186  & !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1  & 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10__dup_186  & (!\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1 
// ))

	.dataa(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_10__dup_186 ),
	.datab(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx44952z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X51_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_11_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_  & \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_  & 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx46946z1  & (!\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_ ))

	.dataa(\u_fir|tap_array_11_filter_block_next_sum_add16_0|nx46946z1 ),
	.datab(\u_fir|tap_array_12_filter_block_prod_mults28_0|d_12_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_12_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X49_Y11_N25
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__15_ ));

// atom is at LCFF_X54_Y11_N17
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__9_ ));

// atom is at LCFF_X49_Y11_N23
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__9_ ));

// atom is at LCFF_X49_Y11_N17
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__8_ ));

// atom is at LCFF_X49_Y11_N19
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__7_ ));

// atom is at LCFF_X54_Y11_N7
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__4_ ));

// atom is at LCFF_X49_Y11_N9
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__4_ ));

// atom is at LCFF_X49_Y11_N15
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__5_ ));

// atom is at LCFF_X54_Y11_N3
cycloneii_lcell_ff \u_fir|tap_array_12_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_11__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_12__2_ ));

// atom is at LCFF_X49_Y11_N5
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__2_ ));

// atom is at LCFF_X49_Y11_N7
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__1_ ));

// atom is at LCCOMB_X49_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52936 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z13  = CARRY(\u_fir|taps_13__0_  & \u_fir|taps_13__2_ )

	.dataa(\u_fir|taps_13__0_ ),
	.datab(\u_fir|taps_13__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52935 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z12  = CARRY(\u_fir|taps_13__3_  & !\u_fir|taps_13__1_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_13__3_  & 
// (!\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_13__1_ ))

	.dataa(\u_fir|taps_13__3_ ),
	.datab(\u_fir|taps_13__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z13 ),
	.combout(),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52934 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11  = CARRY(\u_fir|taps_13__4_  & (\u_fir|taps_13__2_  # !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z12 ) # !\u_fir|taps_13__4_  & \u_fir|taps_13__2_  & 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z12 )

	.dataa(\u_fir|taps_13__4_ ),
	.datab(\u_fir|taps_13__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z12 ),
	.combout(),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52931 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_13__5_  & (\u_fir|taps_13__7_  & \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9  & VCC # !\u_fir|taps_13__7_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9 ) # 
// !\u_fir|taps_13__5_  & (\u_fir|taps_13__7_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_13__7_  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9  # GND))
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z8  = CARRY(\u_fir|taps_13__5_  & !\u_fir|taps_13__7_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9  # !\u_fir|taps_13__5_  & (!\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9  
// # !\u_fir|taps_13__7_ ))

	.dataa(\u_fir|taps_13__5_ ),
	.datab(\u_fir|taps_13__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z9 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52930 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_13__6_  $ \u_fir|taps_13__8_  $ !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z8 ) # GND
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7  = CARRY(\u_fir|taps_13__6_  & (\u_fir|taps_13__8_  # !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z8 ) # !\u_fir|taps_13__6_  & \u_fir|taps_13__8_  & 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z8 )

	.dataa(\u_fir|taps_13__6_ ),
	.datab(\u_fir|taps_13__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z8 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52927 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_13__15_  & (\u_fir|taps_13__9_  & \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5  & VCC # !\u_fir|taps_13__9_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5 ) # 
// !\u_fir|taps_13__15_  & (\u_fir|taps_13__9_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_13__9_  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5  # GND))
// \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z4  = CARRY(\u_fir|taps_13__15_  & !\u_fir|taps_13__9_  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_13__15_  & (!\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5 
//  # !\u_fir|taps_13__9_ ))

	.dataa(\u_fir|taps_13__15_ ),
	.datab(\u_fir|taps_13__9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z5 ),
	.combout(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_prod_mults28_0|modgen_add_13_ix9228z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_  & \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_  & 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx40964z1  & (!\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_ ))

	.dataa(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx40964z1 ),
	.datab(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_13_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_13_filter_block_prod_mults28_0|d_8_  & (!\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_8_ ),
	.datab(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx43955z1  $ \u_fir|tap_array_13_filter_block_prod_mults28_0|d_9_  $ !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx43955z1  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|d_9_  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx43955z1  & \u_fir|tap_array_13_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx43955z1 ),
	.datab(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_13_filter_block_prod_mults28_0|d_11_  $ !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_13_filter_block_prod_mults28_0|d_11_  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_13_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_13_filter_block_prod_mults28_0|d_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z1  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z1  & !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22  
// # !\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z1  & (!\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|tap_array_13_filter_block_prod_mults28_0|nx9228z1 ),
	.datab(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X49_Y11_N21
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__10_ ));

// atom is at LCFF_X46_Y11_N15
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__10_ ));

// atom is at LCFF_X46_Y11_N9
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__7_ ));

// atom is at LCFF_X46_Y11_N5
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__5_ ));

// atom is at LCFF_X46_Y11_N3
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__4_ ));

// atom is at LCFF_X49_Y11_N11
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__3_ ));

// atom is at LCFF_X46_Y11_N1
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__3_ ));

// atom is at LCCOMB_X46_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52939 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx37973z1  = \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx37973z1  & (\u_fir|taps_14__3_  $ VCC) # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|taps_14__3_  & VCC
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46  = CARRY(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx37973z1  & \u_fir|taps_14__3_ )

	.dataa(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx37973z1 ),
	.datab(\u_fir|taps_14__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx37973z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z46 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52939 .lut_mask = 16'h6688;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N4
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|taps_14__5_  $ !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|taps_14__5_  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|taps_14__5_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|taps_14__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N8
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52935 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx41961z1  = (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx41961z1  $ \u_fir|taps_14__7_  $ !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z37 ) # GND
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34  = CARRY(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx41961z1  & (\u_fir|taps_14__7_  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z37 ) # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx41961z1  & \u_fir|taps_14__7_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z37 )

	.dataa(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx41961z1 ),
	.datab(\u_fir|taps_14__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z37 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx41961z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52935 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|taps_14__8_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|taps_14__8_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|taps_14__8_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|taps_14__8_  & 
// (!\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|taps_14__8_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|taps_14__9_  $ \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|taps_14__9_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx43955z1  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z31 ) # !\u_fir|taps_14__9_  & 
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|taps_14__9_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|taps_14__10_  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28  & VCC # !\u_fir|taps_14__10_  & 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|taps_14__10_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|taps_14__10_  & 
// (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|taps_14__10_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx44952z1  & (!\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|taps_14__10_ ))

	.dataa(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx44952z1 ),
	.datab(\u_fir|taps_14__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|taps_14__15_  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|taps_14__15_  & 
// (!\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|taps_14__15_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X46_Y11_N17
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__15_ ));

// atom is at LCFF_X44_Y11_N5
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__15_ ));

// atom is at LCFF_X46_Y11_N13
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__9_ ));

// atom is at LCFF_X44_Y11_N1
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_9_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__9_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__9_ ));

// atom is at LCFF_X44_Y11_N3
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__7_ ));

// atom is at LCFF_X46_Y11_N11
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__8_ ));

// atom is at LCFF_X44_Y12_N31
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__8_ ));

// atom is at LCFF_X44_Y12_N29
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__4_ ));

// atom is at LCFF_X49_Y11_N13
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__6_ ));

// atom is at LCFF_X46_Y11_N7
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__6_ ));

// atom is at LCFF_X44_Y12_N27
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__6_ ));

// atom is at LCFF_X49_Y11_N1
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_13__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__2_ ));

// atom is at LCFF_X44_Y12_N19
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__2_ ));

// atom is at LCCOMB_X49_Y11_N2
cycloneii_lcell_comb \u_fir|taps_14__1_~feeder (
// Equation(s):
// \u_fir|taps_14__1_~feeder_combout  = \u_fir|taps_13__1_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_13__1_ ),
	.cin(gnd),
	.combout(\u_fir|taps_14__1_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_14__1_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_14__1_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X49_Y11_N3
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_14__1_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__1_ ));

// atom is at LCFF_X44_Y12_N23
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__1_ ));

// atom is at LCFF_X44_Y12_N21
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__3_ ));

// atom is at LCCOMB_X44_Y12_N16
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52940 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z17  = CARRY(!\u_fir|taps_15__0_  & !\u_fir|taps_15__1_ )

	.dataa(\u_fir|taps_15__0_ ),
	.datab(\u_fir|taps_15__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z17 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52940 .lut_mask = 16'h0011;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52940 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X44_Y12_N18
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52939 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z16  = CARRY(\u_fir|taps_15__2_  # !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z17 )

	.dataa(vcc),
	.datab(\u_fir|taps_15__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z17 ),
	.combout(),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52939 .lut_mask = 16'h00CF;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52939 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y12_N20
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52938 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z15  = CARRY(\u_fir|taps_15__0_  & (!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z16  # !\u_fir|taps_15__3_ ) # !\u_fir|taps_15__0_  & !\u_fir|taps_15__3_  & 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z16 )

	.dataa(\u_fir|taps_15__0_ ),
	.datab(\u_fir|taps_15__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z16 ),
	.combout(),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z15 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52938 .lut_mask = 16'h002B;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y12_N22
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52937 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z14  = CARRY(\u_fir|taps_15__4_  & (!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z15  # !\u_fir|taps_15__1_ ) # !\u_fir|taps_15__4_  & !\u_fir|taps_15__1_  & 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z15 )

	.dataa(\u_fir|taps_15__4_ ),
	.datab(\u_fir|taps_15__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z15 ),
	.combout(),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z14 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52937 .lut_mask = 16'h002B;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y12_N24
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52936 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13  = CARRY(\u_fir|taps_15__5_  & \u_fir|taps_15__2_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z14  # !\u_fir|taps_15__5_  & (\u_fir|taps_15__2_  # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z14 ))

	.dataa(\u_fir|taps_15__5_ ),
	.datab(\u_fir|taps_15__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z14 ),
	.combout(),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52936 .lut_mask = 16'h004D;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y12_N28
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52934 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_15__7_  $ \u_fir|taps_15__4_  $ \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z12 ) # GND
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11  = CARRY(\u_fir|taps_15__7_  & \u_fir|taps_15__4_  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z12  # !\u_fir|taps_15__7_  & (\u_fir|taps_15__4_  # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z12 ))

	.dataa(\u_fir|taps_15__7_ ),
	.datab(\u_fir|taps_15__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z12 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52934 .lut_mask = 16'h964D;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N0
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52932 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_15__6_  $ \u_fir|taps_15__9_  $ \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z10 ) # GND
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9  = CARRY(\u_fir|taps_15__6_  & (!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z10  # !\u_fir|taps_15__9_ ) # !\u_fir|taps_15__6_  & !\u_fir|taps_15__9_  & 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z10 )

	.dataa(\u_fir|taps_15__6_ ),
	.datab(\u_fir|taps_15__9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z10 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52932 .lut_mask = 16'h962B;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52927 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|d_13_  = !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z5 
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z4  = CARRY(!\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z5 )

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z5 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_13_ ),
	.cout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52927 .lut_mask = 16'h0F0F;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N6
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_  & \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_  & 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx40964z1  & (!\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_ ))

	.dataa(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx40964z1 ),
	.datab(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N12
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_11_  $ \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx43955z1  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_11_  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_11_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_15_filter_block_prod_mults28_0|d_12_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1  & \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_12_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1  & 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_12_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_12_  & (!\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1 ))

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_12_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx44952z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_15_filter_block_prod_mults28_0|d_14_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_14_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_14_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_14_  & (!\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_14_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X44_Y11_N9
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__10_ ));

// atom is at LCFF_X44_Y14_N19
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__10_ ));

// atom is at LCFF_X44_Y14_N15
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__8_ ));

// atom is at LCFF_X44_Y14_N13
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_7_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__7_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__7_ ));

// atom is at LCFF_X44_Y12_N25
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__5_ ));

// atom is at LCFF_X44_Y14_N9
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_5_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__5_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__5_ ));

// atom is at LCFF_X44_Y14_N5
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_3_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__3_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__3_ ));

// atom is at LCFF_X44_Y14_N1
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__1_ ));

// atom is at LCCOMB_X44_Y14_N0
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52936 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z13  = CARRY(\u_fir|taps_16__0_  & \u_fir|taps_16__1_ )

	.dataa(\u_fir|taps_16__0_ ),
	.datab(\u_fir|taps_16__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N2
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52935 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z12  = CARRY(\u_fir|taps_16__2_  & !\u_fir|taps_16__1_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z13  # !\u_fir|taps_16__2_  & 
// (!\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z13  # !\u_fir|taps_16__1_ ))

	.dataa(\u_fir|taps_16__2_ ),
	.datab(\u_fir|taps_16__1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z13 ),
	.combout(),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N4
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52934 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z11  = CARRY(\u_fir|taps_16__2_  & (\u_fir|taps_16__3_  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z12 ) # !\u_fir|taps_16__2_  & \u_fir|taps_16__3_  & 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z12 )

	.dataa(\u_fir|taps_16__2_ ),
	.datab(\u_fir|taps_16__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z12 ),
	.combout(),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N6
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52933 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z10  = CARRY(\u_fir|taps_16__4_  & !\u_fir|taps_16__3_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z11  # !\u_fir|taps_16__4_  & 
// (!\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z11  # !\u_fir|taps_16__3_ ))

	.dataa(\u_fir|taps_16__4_ ),
	.datab(\u_fir|taps_16__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z11 ),
	.combout(),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52933 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N8
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52932 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_16__4_  $ \u_fir|taps_16__5_  $ !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z10 ) # GND
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9  = CARRY(\u_fir|taps_16__4_  & (\u_fir|taps_16__5_  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z10 ) # !\u_fir|taps_16__4_  & \u_fir|taps_16__5_  & 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z10 )

	.dataa(\u_fir|taps_16__4_ ),
	.datab(\u_fir|taps_16__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z10 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N10
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52931 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_16__6_  & (\u_fir|taps_16__5_  & \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9  & VCC # !\u_fir|taps_16__5_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9 ) # 
// !\u_fir|taps_16__6_  & (\u_fir|taps_16__5_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9  # !\u_fir|taps_16__5_  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9  # GND))
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z8  = CARRY(\u_fir|taps_16__6_  & !\u_fir|taps_16__5_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9  # !\u_fir|taps_16__6_  & (!\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9  
// # !\u_fir|taps_16__5_ ))

	.dataa(\u_fir|taps_16__6_ ),
	.datab(\u_fir|taps_16__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z9 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N12
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52930 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_16__6_  $ \u_fir|taps_16__7_  $ !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z8 ) # GND
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7  = CARRY(\u_fir|taps_16__6_  & (\u_fir|taps_16__7_  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z8 ) # !\u_fir|taps_16__6_  & \u_fir|taps_16__7_  & 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z8 )

	.dataa(\u_fir|taps_16__6_ ),
	.datab(\u_fir|taps_16__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z8 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N16
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52928 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_16__9_  $ \u_fir|taps_16__8_  $ !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z6 ) # GND
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5  = CARRY(\u_fir|taps_16__9_  & (\u_fir|taps_16__8_  # !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z6 ) # !\u_fir|taps_16__9_  & \u_fir|taps_16__8_  & 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z6 )

	.dataa(\u_fir|taps_16__9_ ),
	.datab(\u_fir|taps_16__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z6 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N18
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52927 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_16__9_  & (\u_fir|taps_16__10_  & \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5  & VCC # !\u_fir|taps_16__10_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5 ) # 
// !\u_fir|taps_16__9_  & (\u_fir|taps_16__10_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5  # !\u_fir|taps_16__10_  & (\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5  # GND))
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z4  = CARRY(\u_fir|taps_16__9_  & !\u_fir|taps_16__10_  & !\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5  # !\u_fir|taps_16__9_  & (!\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5  
// # !\u_fir|taps_16__10_ ))

	.dataa(\u_fir|taps_16__9_ ),
	.datab(\u_fir|taps_16__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z5 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|modgen_add_15_ix8231z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X44_Y14_N24
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_prod_mults28_0|ix8231z52923 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z1  = \u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z2 ),
	.combout(\u_fir|tap_array_16_filter_block_prod_mults28_0|nx8231z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|ix8231z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_16_filter_block_prod_mults28_0|ix8231z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N6
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_16_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_7_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1  & 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_7_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_7_  & (!\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1 ))

	.dataa(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_7_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx40964z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N14
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_16_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_11_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1  & 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_16_filter_block_prod_mults28_0|d_11_  & (!\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1 ))

	.dataa(\u_fir|tap_array_16_filter_block_prod_mults28_0|d_11_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx44952z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N18
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|taps_16__15_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|taps_16__15_  & 
// (!\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|taps_16__15_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X43_Y14_N23
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_10_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__10_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_10_ ));

// atom is at LCFF_X44_Y14_N21
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__15_ ));

// atom is at LCFF_X43_Y14_N25
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_15_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__15_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_15_ ));

// atom is at LCFF_X43_Y14_N19
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_8_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__8_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_8_ ));

// atom is at LCFF_X44_Y14_N11
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__6_ ));

// atom is at LCFF_X43_Y14_N15
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_6_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__6_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_6_ ));

// atom is at LCFF_X44_Y14_N7
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__4_ ));

// atom is at LCFF_X43_Y14_N11
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_4_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__4_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_4_ ));

// atom is at LCFF_X44_Y14_N3
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__2_ ));

// atom is at LCFF_X43_Y14_N7
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_2_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__2_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_2_ ));

// atom is at LCFF_X43_Y14_N5
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_1_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__1_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_1_ ));

// atom is at LCFF_X53_Y11_N1
cycloneii_lcell_ff \u_fir|tap_array_13_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_12__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_13__0_ ));

// atom is at LCCOMB_X53_Y11_N2
cycloneii_lcell_comb \u_fir|taps_14__0_~feeder (
// Equation(s):
// \u_fir|taps_14__0_~feeder_combout  = \u_fir|taps_13__0_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_fir|taps_13__0_ ),
	.cin(gnd),
	.combout(\u_fir|taps_14__0_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \u_fir|taps_14__0_~feeder .lut_mask = 16'hFF00;
defparam \u_fir|taps_14__0_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X53_Y11_N3
cycloneii_lcell_ff \u_fir|tap_array_14_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\u_fir|taps_14__0_~feeder_combout ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_14__0_ ));

// atom is at LCFF_X44_Y12_N17
cycloneii_lcell_ff \u_fir|tap_array_15_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_14__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_15__0_ ));

// atom is at LCFF_X44_Y12_N9
cycloneii_lcell_ff \u_fir|tap_array_16_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_15__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|taps_16__0_ ));

// atom is at LCFF_X43_Y14_N3
cycloneii_lcell_ff \u_fir|tap_array_17_filter_block_reg_current_tap_0_ (
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(gnd),
	.sdata(\u_fir|taps_16__0_ ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_fir|tap_array_17_filter_block_tap_next_0_ ));

// atom is at LCCOMB_X43_Y14_N2
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52938 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z15  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_3_  & \u_fir|tap_array_17_filter_block_tap_next_0_ )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_3_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_0_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z15 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52938 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52938 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N4
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52937 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z14  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_4_  & !\u_fir|tap_array_17_filter_block_tap_next_1_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z15  # 
// !\u_fir|tap_array_17_filter_block_tap_next_4_  & (!\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z15  # !\u_fir|tap_array_17_filter_block_tap_next_1_ ))

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_4_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z15 ),
	.combout(),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z14 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52937 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N6
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52936 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_5_  & (\u_fir|tap_array_17_filter_block_tap_next_2_  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z14 ) # 
// !\u_fir|tap_array_17_filter_block_tap_next_5_  & \u_fir|tap_array_17_filter_block_tap_next_2_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z14 )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_5_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z14 ),
	.combout(),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52936 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N8
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52935 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_3_  = \u_fir|tap_array_17_filter_block_tap_next_3_  & (\u_fir|tap_array_17_filter_block_tap_next_6_  & \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13  & VCC # 
// !\u_fir|tap_array_17_filter_block_tap_next_6_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13 ) # !\u_fir|tap_array_17_filter_block_tap_next_3_  & (\u_fir|tap_array_17_filter_block_tap_next_6_  & 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13  # !\u_fir|tap_array_17_filter_block_tap_next_6_  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13  # GND))
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z12  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_3_  & !\u_fir|tap_array_17_filter_block_tap_next_6_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13  # 
// !\u_fir|tap_array_17_filter_block_tap_next_3_  & (!\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13  # !\u_fir|tap_array_17_filter_block_tap_next_6_ ))

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_3_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z13 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52935 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N10
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52934 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_  = (\u_fir|tap_array_17_filter_block_tap_next_7_  $ \u_fir|tap_array_17_filter_block_tap_next_4_  $ !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z12 ) # GND
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_7_  & (\u_fir|tap_array_17_filter_block_tap_next_4_  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z12 ) # 
// !\u_fir|tap_array_17_filter_block_tap_next_7_  & \u_fir|tap_array_17_filter_block_tap_next_4_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z12 )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_7_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z12 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52934 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N12
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52933 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_5_  = \u_fir|tap_array_17_filter_block_tap_next_5_  & (\u_fir|tap_array_17_filter_block_tap_next_8_  & \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11  & VCC # 
// !\u_fir|tap_array_17_filter_block_tap_next_8_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11 ) # !\u_fir|tap_array_17_filter_block_tap_next_5_  & (\u_fir|tap_array_17_filter_block_tap_next_8_  & 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11  # !\u_fir|tap_array_17_filter_block_tap_next_8_  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11  # GND))
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z10  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_5_  & !\u_fir|tap_array_17_filter_block_tap_next_8_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11  # 
// !\u_fir|tap_array_17_filter_block_tap_next_5_  & (!\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11  # !\u_fir|tap_array_17_filter_block_tap_next_8_ ))

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_5_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z11 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N16
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52931 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_7_  = \u_fir|tap_array_17_filter_block_tap_next_7_  & (\u_fir|tap_array_17_filter_block_tap_next_10_  & \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9  & VCC # 
// !\u_fir|tap_array_17_filter_block_tap_next_10_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9 ) # !\u_fir|tap_array_17_filter_block_tap_next_7_  & (\u_fir|tap_array_17_filter_block_tap_next_10_  & 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9  # !\u_fir|tap_array_17_filter_block_tap_next_10_  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9  # GND))
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z8  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_7_  & !\u_fir|tap_array_17_filter_block_tap_next_10_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9  # 
// !\u_fir|tap_array_17_filter_block_tap_next_7_  & (!\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9  # !\u_fir|tap_array_17_filter_block_tap_next_10_ ))

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_7_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z9 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52931 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N18
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52930 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_  = (\u_fir|tap_array_17_filter_block_tap_next_15_  $ \u_fir|tap_array_17_filter_block_tap_next_8_  $ !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z8 ) # GND
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_15_  & (\u_fir|tap_array_17_filter_block_tap_next_8_  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z8 ) # 
// !\u_fir|tap_array_17_filter_block_tap_next_15_  & \u_fir|tap_array_17_filter_block_tap_next_8_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z8 )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z8 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N20
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52929 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_9_  = \u_fir|tap_array_17_filter_block_tap_next_9_  & (\u_fir|tap_array_17_filter_block_tap_next_15_  & \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7  & VCC # 
// !\u_fir|tap_array_17_filter_block_tap_next_15_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7 ) # !\u_fir|tap_array_17_filter_block_tap_next_9_  & (\u_fir|tap_array_17_filter_block_tap_next_15_  & 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7  # !\u_fir|tap_array_17_filter_block_tap_next_15_  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7  # GND))
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z6  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_9_  & !\u_fir|tap_array_17_filter_block_tap_next_15_  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7  # 
// !\u_fir|tap_array_17_filter_block_tap_next_9_  & (!\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7  # !\u_fir|tap_array_17_filter_block_tap_next_15_ ))

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_9_ ),
	.datab(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z7 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X43_Y14_N24
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52927 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_prod_mults28_0|d_11_  = (\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z5 ) # GND
// \u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z4  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_15_ )

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z5 ),
	.combout(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_11_ ),
	.cout(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52927 .lut_mask = 16'hF0AA;
defparam \u_fir|tap_array_17_filter_block_prod_mults28_0|ix12219z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N4
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|tap_array_17_filter_block_prod_mults28_0|d_5_  $ !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_5_  # !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|tap_array_17_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N6
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_17_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1  & \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1  & 
// !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_6_  & (!\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1 ))

	.dataa(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_6_ ),
	.datab(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx40964z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N12
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx43955z1  $ \u_fir|tap_array_17_filter_block_prod_mults28_0|d_9_  $ !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx43955z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_9_  # !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx43955z1  & \u_fir|tap_array_17_filter_block_prod_mults28_0|d_9_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx43955z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N14
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_17_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1  & \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1  & 
// !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_10_  & (!\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1 ))

	.dataa(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx44952z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N16
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52931 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx45949z1  = (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx45949z1  $ \u_fir|tap_array_17_filter_block_prod_mults28_0|d_11_  $ !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z25 ) # GND
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx45949z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_11_  # !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z25 ) # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx45949z1  & \u_fir|tap_array_17_filter_block_prod_mults28_0|d_11_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z25 )

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx45949z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z25 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx45949z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52931 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N18
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52930 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx46946z1  = \u_fir|tap_array_17_filter_block_prod_mults28_0|d_12_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1  & \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22  & VCC # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22 ) # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_12_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1  & 
// !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1  & (\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22  # GND))
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z19  = CARRY(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_12_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22  # 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_12_  & (!\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1 ))

	.dataa(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_12_ ),
	.datab(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx46946z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z22 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx46946z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52930 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at PIN_V1
cycloneii_io sw_ibuf_16_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(\sw~combout [16]),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[16]));
// synopsys translate_off
defparam sw_ibuf_16_.input_async_reset = "none";
defparam sw_ibuf_16_.input_power_up = "low";
defparam sw_ibuf_16_.input_register_mode = "none";
defparam sw_ibuf_16_.input_sync_reset = "none";
defparam sw_ibuf_16_.oe_async_reset = "none";
defparam sw_ibuf_16_.oe_power_up = "low";
defparam sw_ibuf_16_.oe_register_mode = "none";
defparam sw_ibuf_16_.oe_sync_reset = "none";
defparam sw_ibuf_16_.operation_mode = "input";
defparam sw_ibuf_16_.output_async_reset = "none";
defparam sw_ibuf_16_.output_power_up = "low";
defparam sw_ibuf_16_.output_register_mode = "none";
defparam sw_ibuf_16_.output_sync_reset = "none";
// synopsys translate_on

// atom is at LCFF_X34_Y14_N29
cycloneii_lcell_ff reg_audio_out_9_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_9_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx46946z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_9_));

// atom is at LCCOMB_X34_Y14_N30
cycloneii_lcell_comb ix50814z52923(
// Equation(s):
// nx50814z1 = bit_position_1_ $ bit_position_0_

	.dataa(vcc),
	.datab(vcc),
	.datac(bit_position_1_),
	.datad(bit_position_0_),
	.cin(gnd),
	.combout(nx50814z1),
	.cout());
// synopsys translate_off
defparam ix50814z52923.lut_mask = 16'h0FF0;
defparam ix50814z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y14_N31
cycloneii_lcell_ff modgen_counter_bit_position_reg_q_1_(
	.clk(\aud_bclk_dup0~clkctrl_outclk ),
	.datain(nx50814z1),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(bit_position_1_));

// atom is at LCFF_X34_Y14_N23
cycloneii_lcell_ff reg_audio_out_8_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_8_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx45949z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_8_));

// atom is at LCCOMB_X35_Y14_N2
cycloneii_lcell_comb ix24999z52930(
// Equation(s):
// nx24999z7 = bit_position_0_ & (bit_position_1_ & audio_out_8_) # !bit_position_0_ & (audio_out_9_ # !bit_position_1_)

	.dataa(bit_position_0_),
	.datab(audio_out_9_),
	.datac(bit_position_1_),
	.datad(audio_out_8_),
	.cin(gnd),
	.combout(nx24999z7),
	.cout());
// synopsys translate_off
defparam ix24999z52930.lut_mask = 16'hE545;
defparam ix24999z52930.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N20
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx62798z1  $ \u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  $ !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx62798z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  # !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx62798z1  & \u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx62798z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X35_Y14_N21
cycloneii_lcell_ff reg_audio_out_10_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_10_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx62798z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_10_));

// atom is at LCCOMB_X42_Y14_N22
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  & \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  & 
// !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  & (\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx63795z1  & (!\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_ ))

	.dataa(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx63795z1 ),
	.datab(\u_fir|tap_array_17_filter_block_prod_mults28_0|d_13_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X35_Y14_N15
cycloneii_lcell_ff reg_audio_out_11_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_11_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx63795z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_11_));

// atom is at LCCOMB_X35_Y14_N8
cycloneii_lcell_comb ix24999z52929(
// Equation(s):
// nx24999z6 = bit_position_1_ & nx24999z7 # !bit_position_1_ & (nx24999z7 & (audio_out_11_) # !nx24999z7 & audio_out_10_)

	.dataa(bit_position_1_),
	.datab(nx24999z7),
	.datac(audio_out_10_),
	.datad(audio_out_11_),
	.cin(gnd),
	.combout(nx24999z6),
	.cout());
// synopsys translate_off
defparam ix24999z52929.lut_mask = 16'hDC98;
defparam ix24999z52929.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y14_N19
cycloneii_lcell_ff reg_audio_out_7_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_7_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx44952z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_7_));

// atom is at LCFF_X34_Y14_N17
cycloneii_lcell_ff reg_audio_out_6_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_6_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx43955z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_6_));

// atom is at LCCOMB_X35_Y14_N26
cycloneii_lcell_comb ix24999z52925(
// Equation(s):
// nx24999z2 = nx24999z3 & (audio_out_7_ # bit_position_1_) # !nx24999z3 & (!bit_position_1_ & audio_out_6_)

	.dataa(nx24999z3),
	.datab(audio_out_7_),
	.datac(bit_position_1_),
	.datad(audio_out_6_),
	.cin(gnd),
	.combout(nx24999z2),
	.cout());
// synopsys translate_off
defparam ix24999z52925.lut_mask = 16'hADA8;
defparam ix24999z52925.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X31_Y14_N23
cycloneii_lcell_ff reg_audio_out_3_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_3_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx40964z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_3_));

// atom is at LCFF_X34_Y14_N11
cycloneii_lcell_ff reg_audio_out_2_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(raw_audio_2_),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx39967z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_2_));

// atom is at LCCOMB_X35_Y14_N4
cycloneii_lcell_comb ix24999z52927(
// Equation(s):
// nx24999z4 = nx24999z5 & (audio_out_3_ # bit_position_1_) # !nx24999z5 & (!bit_position_1_ & audio_out_2_)

	.dataa(nx24999z5),
	.datab(audio_out_3_),
	.datac(bit_position_1_),
	.datad(audio_out_2_),
	.cin(gnd),
	.combout(nx24999z4),
	.cout());
// synopsys translate_off
defparam ix24999z52927.lut_mask = 16'hADA8;
defparam ix24999z52927.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X35_Y14_N24
cycloneii_lcell_comb ix24999z52924(
// Equation(s):
// nx24999z1 = bit_position_3_ & (bit_position_2_ & (nx24999z4) # !bit_position_2_ & nx24999z2) # !bit_position_3_ & (!bit_position_2_)

	.dataa(bit_position_3_),
	.datab(nx24999z2),
	.datac(nx24999z4),
	.datad(bit_position_2_),
	.cin(gnd),
	.combout(nx24999z1),
	.cout());
// synopsys translate_off
defparam ix24999z52924.lut_mask = 16'hA0DD;
defparam ix24999z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X35_Y14_N18
cycloneii_lcell_comb \audio_out_13_~feeder (
// Equation(s):
// \audio_out_13_~feeder_combout  = raw_audio_11_

	.dataa(vcc),
	.datab(raw_audio_11_),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\audio_out_13_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \audio_out_13_~feeder .lut_mask = 16'hCCCC;
defparam \audio_out_13_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X44_Y11_N16
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52923 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  = \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z2 ),
	.combout(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_15_filter_block_prod_mults28_0|ix15210z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52927 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_9__9_  & (\u_fir|taps_9__10_  & \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5  & VCC # !\u_fir|taps_9__10_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5 ) # 
// !\u_fir|taps_9__9_  & (\u_fir|taps_9__10_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_9__10_  & (\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5  # GND))
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z4  = CARRY(\u_fir|taps_9__9_  & !\u_fir|taps_9__10_  & !\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_9__9_  & (!\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5  # 
// !\u_fir|taps_9__10_ ))

	.dataa(\u_fir|taps_9__9_ ),
	.datab(\u_fir|taps_9__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z5 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|modgen_add_8_ix9228z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y11_N28
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_prod_mults28_0|ix9228z52923 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1  = \u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z2 ),
	.combout(\u_fir|tap_array_9_filter_block_prod_mults28_0|nx9228z1 ),
	.cout());
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|ix9228z52923 .lut_mask = 16'hF0F0;
defparam \u_fir|tap_array_9_filter_block_prod_mults28_0|ix9228z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N16
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52932 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_6__9_  $ \u_fir|taps_6__8_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z9 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8  = CARRY(\u_fir|taps_6__9_  & (\u_fir|taps_6__8_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z9 ) # !\u_fir|taps_6__9_  & \u_fir|taps_6__8_  & 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z9 )

	.dataa(\u_fir|taps_6__9_ ),
	.datab(\u_fir|taps_6__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z9 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z8 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52932 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y9_N20
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52930 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_10_  = (\u_fir|taps_6__15_  $ \u_fir|taps_6__10_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z7 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z6  = CARRY(\u_fir|taps_6__15_  & (\u_fir|taps_6__10_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z7 ) # !\u_fir|taps_6__15_  & \u_fir|taps_6__10_  & 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z7 )

	.dataa(\u_fir|taps_6__15_ ),
	.datab(\u_fir|taps_6__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z7 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10_ ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_4_ix10225z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N14
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52943 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_7__dup_189  = \u_fir|tap_array_6_filter_block_prod_mults28_0|d_9_  & (\u_fir|taps_6__7_  & \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20  & VCC # !\u_fir|taps_6__7_  & 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20 ) # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9_  & (\u_fir|taps_6__7_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20  # !\u_fir|taps_6__7_  & 
// (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20  # GND))
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z19  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9_  & !\u_fir|taps_6__7_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20  # 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9_  & (!\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20  # !\u_fir|taps_6__7_ ))

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9_ ),
	.datab(\u_fir|taps_6__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z20 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_7__dup_189 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z19 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52943 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52943 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y9_N20
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52927 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186  = (\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z5  $ \u_fir|taps_6__10_  $ !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z17 ) # GND
// \u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z4  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z5  & (\u_fir|taps_6__10_  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z17 ) # 
// !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z5  & \u_fir|taps_6__10_  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z17 )

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z5 ),
	.datab(\u_fir|taps_6__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z17 ),
	.combout(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186 ),
	.cout(\u_fir|tap_array_6_filter_block_prod_mults28_0|nx10225z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_prod_mults28_0|modgen_add_5_ix10225z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N4
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52936 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z13  = CARRY(\u_fir|taps_5__0_  & \u_fir|taps_5__2_ )

	.dataa(\u_fir|taps_5__0_ ),
	.datab(\u_fir|taps_5__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N6
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52935 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z12  = CARRY(\u_fir|taps_5__1_  & !\u_fir|taps_5__3_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z13  # !\u_fir|taps_5__1_  & (!\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z13  # 
// !\u_fir|taps_5__3_ ))

	.dataa(\u_fir|taps_5__1_ ),
	.datab(\u_fir|taps_5__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z13 ),
	.combout(),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N8
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52934 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11  = CARRY(\u_fir|taps_5__2_  & (\u_fir|taps_5__4_  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z12 ) # !\u_fir|taps_5__2_  & \u_fir|taps_5__4_  & 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z12 )

	.dataa(\u_fir|taps_5__2_ ),
	.datab(\u_fir|taps_5__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z12 ),
	.combout(),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N16
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52930 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_5__6_  $ \u_fir|taps_5__8_  $ !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z8 ) # GND
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7  = CARRY(\u_fir|taps_5__6_  & (\u_fir|taps_5__8_  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z8 ) # !\u_fir|taps_5__6_  & \u_fir|taps_5__8_  & 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z8 )

	.dataa(\u_fir|taps_5__6_ ),
	.datab(\u_fir|taps_5__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z8 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52930 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X55_Y12_N18
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52929 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_5__9_  & (\u_fir|taps_5__7_  & \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7  & VCC # !\u_fir|taps_5__7_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7 ) # 
// !\u_fir|taps_5__9_  & (\u_fir|taps_5__7_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_5__7_  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7  # GND))
// \u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z6  = CARRY(\u_fir|taps_5__9_  & !\u_fir|taps_5__7_  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_5__9_  & (!\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7  # 
// !\u_fir|taps_5__7_ ))

	.dataa(\u_fir|taps_5__9_ ),
	.datab(\u_fir|taps_5__7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z7 ),
	.combout(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_5_filter_block_prod_mults28_0|nx9228z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_prod_mults28_0|modgen_add_3_ix9228z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N0
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52936 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z13  = CARRY(\u_fir|taps_2__1_  & \u_fir|taps_2__0_ )

	.dataa(\u_fir|taps_2__1_ ),
	.datab(\u_fir|taps_2__0_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52936 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N2
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52935 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z12  = CARRY(\u_fir|taps_2__1_  & !\u_fir|taps_2__2_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z13  # !\u_fir|taps_2__1_  & (!\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z13  # 
// !\u_fir|taps_2__2_ ))

	.dataa(\u_fir|taps_2__1_ ),
	.datab(\u_fir|taps_2__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z13 ),
	.combout(),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52935 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N4
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52934 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z11  = CARRY(\u_fir|taps_2__3_  & (\u_fir|taps_2__2_  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z12 ) # !\u_fir|taps_2__3_  & \u_fir|taps_2__2_  & 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z12 )

	.dataa(\u_fir|taps_2__3_ ),
	.datab(\u_fir|taps_2__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z12 ),
	.combout(),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52934 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N6
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52933 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z10  = CARRY(\u_fir|taps_2__4_  & !\u_fir|taps_2__3_  & !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z11  # !\u_fir|taps_2__4_  & (!\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z11  # 
// !\u_fir|taps_2__3_ ))

	.dataa(\u_fir|taps_2__4_ ),
	.datab(\u_fir|taps_2__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z11 ),
	.combout(),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52933 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X49_Y16_N16
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52928 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_2__9_  $ \u_fir|taps_2__8_  $ !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z6 ) # GND
// \u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5  = CARRY(\u_fir|taps_2__9_  & (\u_fir|taps_2__8_  # !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z6 ) # !\u_fir|taps_2__9_  & \u_fir|taps_2__8_  & 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z6 )

	.dataa(\u_fir|taps_2__9_ ),
	.datab(\u_fir|taps_2__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z6 ),
	.combout(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_2_filter_block_prod_mults28_0|nx8231z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_prod_mults28_0|modgen_add_1_ix8231z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N0
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52938 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z15  = CARRY(\u_fir|taps_1__3_  & \u_fir|taps_1__0_ )

	.dataa(\u_fir|taps_1__3_ ),
	.datab(\u_fir|taps_1__0_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z15 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52938 .lut_mask = 16'h0088;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52938 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N2
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52937 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z14  = CARRY(\u_fir|taps_1__1_  & !\u_fir|taps_1__4_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z15  # !\u_fir|taps_1__1_  & (!\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z15  
// # !\u_fir|taps_1__4_ ))

	.dataa(\u_fir|taps_1__1_ ),
	.datab(\u_fir|taps_1__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z15 ),
	.combout(),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z14 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52937 .lut_mask = 16'h0017;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N4
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52936 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13  = CARRY(\u_fir|taps_1__5_  & (\u_fir|taps_1__2_  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z14 ) # !\u_fir|taps_1__5_  & \u_fir|taps_1__2_  & 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z14 )

	.dataa(\u_fir|taps_1__5_ ),
	.datab(\u_fir|taps_1__2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z14 ),
	.combout(),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52936 .lut_mask = 16'h008E;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N6
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52935 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_3_  = \u_fir|taps_1__6_  & (\u_fir|taps_1__3_  & \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13  & VCC # !\u_fir|taps_1__3_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13 ) # 
// !\u_fir|taps_1__6_  & (\u_fir|taps_1__3_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13  # !\u_fir|taps_1__3_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13  # GND))
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z12  = CARRY(\u_fir|taps_1__6_  & !\u_fir|taps_1__3_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13  # !\u_fir|taps_1__6_  & (!\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13  
// # !\u_fir|taps_1__3_ ))

	.dataa(\u_fir|taps_1__6_ ),
	.datab(\u_fir|taps_1__3_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z13 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_3_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52935 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N8
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52934 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_  = (\u_fir|taps_1__7_  $ \u_fir|taps_1__4_  $ !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z12 ) # GND
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11  = CARRY(\u_fir|taps_1__7_  & (\u_fir|taps_1__4_  # !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z12 ) # !\u_fir|taps_1__7_  & \u_fir|taps_1__4_  & 
// !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z12 )

	.dataa(\u_fir|taps_1__7_ ),
	.datab(\u_fir|taps_1__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z12 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_4_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52934 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X48_Y16_N10
cycloneii_lcell_comb \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52933 (
// Equation(s):
// \u_fir|tap_array_1_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_1__5_  & (\u_fir|taps_1__8_  & \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11  & VCC # !\u_fir|taps_1__8_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11 ) # 
// !\u_fir|taps_1__5_  & (\u_fir|taps_1__8_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11  # !\u_fir|taps_1__8_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11  # GND))
// \u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z10  = CARRY(\u_fir|taps_1__5_  & !\u_fir|taps_1__8_  & !\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11  # !\u_fir|taps_1__5_  & (!\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11  
// # !\u_fir|taps_1__8_ ))

	.dataa(\u_fir|taps_1__5_ ),
	.datab(\u_fir|taps_1__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z11 ),
	.combout(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_1_filter_block_prod_mults28_0|nx12219z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52933 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_1_filter_block_prod_mults28_0|ix12219z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y16_N4
cycloneii_lcell_comb \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_2_filter_block_prod_mults28_0|d_6_  $ \u_fir|tap_array_1_filter_block_prod_mults28_0|d_5_  $ !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_1_filter_block_prod_mults28_0|d_5_  # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_2_filter_block_prod_mults28_0|d_6_  & \u_fir|tap_array_1_filter_block_prod_mults28_0|d_5_  & !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_2_filter_block_prod_mults28_0|d_6_ ),
	.datab(\u_fir|tap_array_1_filter_block_prod_mults28_0|d_5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_2_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y16_N16
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52940 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z17  = CARRY(!\u_fir|taps_3__1_  & !\u_fir|taps_3__0_ )

	.dataa(\u_fir|taps_3__1_ ),
	.datab(\u_fir|taps_3__0_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z17 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52940 .lut_mask = 16'h0011;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52940 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X53_Y16_N18
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52939 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z16  = CARRY(\u_fir|taps_3__2_  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z17 )

	.dataa(\u_fir|taps_3__2_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z17 ),
	.combout(),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52939 .lut_mask = 16'h00AF;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52939 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y16_N20
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52938 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z15  = CARRY(\u_fir|taps_3__3_  & \u_fir|taps_3__0_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z16  # !\u_fir|taps_3__3_  & (\u_fir|taps_3__0_  # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z16 ))

	.dataa(\u_fir|taps_3__3_ ),
	.datab(\u_fir|taps_3__0_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z16 ),
	.combout(),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z15 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52938 .lut_mask = 16'h004D;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y16_N22
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52937 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z14  = CARRY(\u_fir|taps_3__1_  & \u_fir|taps_3__4_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z15  # !\u_fir|taps_3__1_  & (\u_fir|taps_3__4_  # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z15 ))

	.dataa(\u_fir|taps_3__1_ ),
	.datab(\u_fir|taps_3__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z15 ),
	.combout(),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z14 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52937 .lut_mask = 16'h004D;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y16_N24
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52936 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13  = CARRY(\u_fir|taps_3__2_  & (!\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z14  # !\u_fir|taps_3__5_ ) # !\u_fir|taps_3__2_  & !\u_fir|taps_3__5_  & 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z14 )

	.dataa(\u_fir|taps_3__2_ ),
	.datab(\u_fir|taps_3__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z14 ),
	.combout(),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52936 .lut_mask = 16'h002B;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y16_N26
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52935 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_5_  = \u_fir|taps_3__3_  & (\u_fir|taps_3__6_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13  # !\u_fir|taps_3__6_  & \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13  & VCC) # 
// !\u_fir|taps_3__3_  & (\u_fir|taps_3__6_  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13  # GND) # !\u_fir|taps_3__6_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13 )
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z12  = CARRY(\u_fir|taps_3__3_  & \u_fir|taps_3__6_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13  # !\u_fir|taps_3__3_  & (\u_fir|taps_3__6_  # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13 ))

	.dataa(\u_fir|taps_3__3_ ),
	.datab(\u_fir|taps_3__6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z13 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_5_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z12 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52935 .lut_mask = 16'h694D;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y16_N28
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52934 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_  = (\u_fir|taps_3__7_  $ \u_fir|taps_3__4_  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z12 ) # GND
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11  = CARRY(\u_fir|taps_3__7_  & \u_fir|taps_3__4_  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z12  # !\u_fir|taps_3__7_  & (\u_fir|taps_3__4_  # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z12 ))

	.dataa(\u_fir|taps_3__7_ ),
	.datab(\u_fir|taps_3__4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z12 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_6_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z11 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52934 .lut_mask = 16'h964D;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X53_Y15_N0
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52932 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_3__6_  $ \u_fir|taps_3__9_  $ \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z10 ) # GND
// \u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9  = CARRY(\u_fir|taps_3__6_  & (!\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z10  # !\u_fir|taps_3__9_ ) # !\u_fir|taps_3__6_  & !\u_fir|taps_3__9_  & 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z10 )

	.dataa(\u_fir|taps_3__6_ ),
	.datab(\u_fir|taps_3__9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z10 ),
	.combout(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_3_filter_block_prod_mults28_0|nx15210z9 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52932 .lut_mask = 16'h962B;
defparam \u_fir|tap_array_3_filter_block_prod_mults28_0|ix15210z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y16_N6
cycloneii_lcell_comb \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_2_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_  & \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_  & 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx40964z1  & (!\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_ ))

	.dataa(\u_fir|tap_array_2_filter_block_next_sum_add16_0|nx40964z1 ),
	.datab(\u_fir|tap_array_3_filter_block_prod_mults28_0|d_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_3_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y12_N4
cycloneii_lcell_comb \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52937 (
// Equation(s):
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx39967z1  = (\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx39967z1  $ \u_fir|taps_4__5_  $ !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z43 ) # GND
// \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40  = CARRY(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx39967z1  & (\u_fir|taps_4__5_  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z43 ) # 
// !\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx39967z1  & \u_fir|taps_4__5_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z43 )

	.dataa(\u_fir|tap_array_3_filter_block_next_sum_add16_0|nx39967z1 ),
	.datab(\u_fir|taps_4__5_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z43 ),
	.combout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx39967z1 ),
	.cout(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx2247z40 ));
// synopsys translate_off
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52937 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_4_filter_block_next_sum_add16_0|ix2247z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N6
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52936 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1  = \u_fir|tap_array_4_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40  & VCC # 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40 ) # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx40964z1  & (\u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_  & 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40  # GND))
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z37  = CARRY(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx40964z1  & !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40  # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx40964z1  & (!\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40  # !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_ ))

	.dataa(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx40964z1 ),
	.datab(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_6_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z40 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx40964z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z37 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52936 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y12_N10
cycloneii_lcell_comb \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_5_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_5_filter_block_prod_mults28_0|d_8_  & (!\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|tap_array_5_filter_block_prod_mults28_0|d_8_ ),
	.datab(\u_fir|tap_array_4_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_5_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N10
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_6_filter_block_prod_mults28_0|d_8__dup_188  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_8__dup_188  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_8__dup_188  & !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34  
// # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_8__dup_188  & (!\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_8__dup_188 ),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N12
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9__dup_187  $ \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9__dup_187  & (\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx43955z1  # !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z31 ) 
// # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9__dup_187  & \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_9__dup_187 ),
	.datab(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y10_N14
cycloneii_lcell_comb \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_5_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28  & VCC 
// # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186 
//  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186  & !\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28  
// # !\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx44952z1  & (!\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186 ))

	.dataa(\u_fir|tap_array_5_filter_block_next_sum_add16_0|nx44952z1 ),
	.datab(\u_fir|tap_array_6_filter_block_prod_mults28_0|d_10__dup_186 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_6_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X58_Y10_N12
cycloneii_lcell_comb \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52933 (
// Equation(s):
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx43955z1  = (\u_fir|tap_array_7_filter_block_prod_mults28_0|d_9_  $ \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx43955z1  $ !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z31 ) # GND
// \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28  = CARRY(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_9_  & (\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx43955z1  # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z31 ) # 
// !\u_fir|tap_array_7_filter_block_prod_mults28_0|d_9_  & \u_fir|tap_array_6_filter_block_next_sum_add16_0|nx43955z1  & !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z31 )

	.dataa(\u_fir|tap_array_7_filter_block_prod_mults28_0|d_9_ ),
	.datab(\u_fir|tap_array_6_filter_block_next_sum_add16_0|nx43955z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z31 ),
	.combout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx43955z1 ),
	.cout(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx2247z28 ));
// synopsys translate_off
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52933 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_7_filter_block_next_sum_add16_0|ix2247z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N18
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52929 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_7_  = \u_fir|taps_8__7_  & (\u_fir|taps_8__8_  & \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7  & VCC # !\u_fir|taps_8__8_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7 ) # 
// !\u_fir|taps_8__7_  & (\u_fir|taps_8__8_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_8__8_  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7  # GND))
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z6  = CARRY(\u_fir|taps_8__7_  & !\u_fir|taps_8__8_  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7  # !\u_fir|taps_8__7_  & (!\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7  # 
// !\u_fir|taps_8__8_ ))

	.dataa(\u_fir|taps_8__7_ ),
	.datab(\u_fir|taps_8__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z7 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_7_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z6 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52929 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y9_N20
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52928 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_  = (\u_fir|taps_8__9_  $ \u_fir|taps_8__8_  $ !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z6 ) # GND
// \u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5  = CARRY(\u_fir|taps_8__9_  & (\u_fir|taps_8__8_  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z6 ) # !\u_fir|taps_8__9_  & \u_fir|taps_8__8_  & 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z6 )

	.dataa(\u_fir|taps_8__9_ ),
	.datab(\u_fir|taps_8__8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z6 ),
	.combout(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_ ),
	.cout(\u_fir|tap_array_8_filter_block_prod_mults28_0|nx9228z5 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52928 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_8_filter_block_prod_mults28_0|modgen_add_7_ix9228z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N10
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_  & 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx42958z1  & (!\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_ ))

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx42958z1 ),
	.datab(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_8_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y10_N14
cycloneii_lcell_comb \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_7_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_  & \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_  & 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx44952z1  & (!\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_ ))

	.dataa(\u_fir|tap_array_7_filter_block_next_sum_add16_0|nx44952z1 ),
	.datab(\u_fir|tap_array_8_filter_block_prod_mults28_0|d_10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_8_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N10
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52934 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1  = \u_fir|tap_array_9_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34  & VCC # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34 ) # !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_8_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1  & 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34  # GND))
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z31  = CARRY(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_8_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34  # 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_8_  & (!\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1 ))

	.dataa(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_8_ ),
	.datab(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx42958z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z34 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx42958z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z31 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52934 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y11_N14
cycloneii_lcell_comb \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52932 (
// Equation(s):
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1  = \u_fir|tap_array_9_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1  & \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28  & VCC # 
// !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28 ) # !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_10_  & (\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1  & 
// !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1  & (\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28  # GND))
// \u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z25  = CARRY(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_10_  & !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1  & !\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28  # 
// !\u_fir|tap_array_9_filter_block_prod_mults28_0|d_10_  & (!\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28  # !\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1 ))

	.dataa(\u_fir|tap_array_9_filter_block_prod_mults28_0|d_10_ ),
	.datab(\u_fir|tap_array_8_filter_block_next_sum_add16_0|nx44952z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z28 ),
	.combout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx44952z1 ),
	.cout(\u_fir|tap_array_9_filter_block_next_sum_add16_0|nx2247z25 ));
// synopsys translate_off
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52932 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_9_filter_block_next_sum_add16_0|ix2247z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X57_Y11_N18
cycloneii_lcell_comb \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52927 (
// Equation(s):
// \u_fir|tap_array_10_filter_block_prod_mults28_0|d_9_  = \u_fir|taps_10__9_  & (\u_fir|taps_10__10_  & \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5  & VCC # !\u_fir|taps_10__10_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5 ) # 
// !\u_fir|taps_10__9_  & (\u_fir|taps_10__10_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_10__10_  & (\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5  # GND))
// \u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z4  = CARRY(\u_fir|taps_10__9_  & !\u_fir|taps_10__10_  & !\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5  # !\u_fir|taps_10__9_  & (!\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5  
// # !\u_fir|taps_10__10_ ))

	.dataa(\u_fir|taps_10__9_ ),
	.datab(\u_fir|taps_10__10_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z5 ),
	.combout(\u_fir|tap_array_10_filter_block_prod_mults28_0|d_9_ ),
	.cout(\u_fir|tap_array_10_filter_block_prod_mults28_0|nx9228z4 ));
// synopsys translate_off
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52927 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_10_filter_block_prod_mults28_0|modgen_add_9_ix9228z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X50_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|taps_13__15_  $ \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx62798z1  $ !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|taps_13__15_  & (\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx62798z1  # !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z19 ) # !\u_fir|taps_13__15_  & 
// \u_fir|tap_array_12_filter_block_next_sum_add16_0|nx62798z1  & !\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|taps_13__15_ ),
	.datab(\u_fir|tap_array_12_filter_block_next_sum_add16_0|nx62798z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_13_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X46_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|taps_14__15_  $ \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx62798z1  $ !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|taps_14__15_  & (\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx62798z1  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z19 ) # !\u_fir|taps_14__15_  & 
// \u_fir|tap_array_13_filter_block_next_sum_add16_0|nx62798z1  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|taps_14__15_ ),
	.datab(\u_fir|tap_array_13_filter_block_next_sum_add16_0|nx62798z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_14_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N20
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52929 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx62798z1  = (\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_  $ \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx62798z1  $ !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z19 ) # GND
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx62798z1  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z19 ) # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_  & \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx62798z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z19 )

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx62798z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z19 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx62798z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52929 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N22
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52928 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1  = \u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1  & \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16  & VCC # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16 ) # !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_  & (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1  & 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16  # GND))
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z13  = CARRY(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_  & !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16  # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_  & (!\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16  # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1 ))

	.dataa(\u_fir|tap_array_15_filter_block_prod_mults28_0|d_15_ ),
	.datab(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx63795z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z16 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx63795z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z13 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52928 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N24
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx64792z1  $ \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  $ !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z13 ) # 
// GND
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx64792z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z13 
// ) # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx64792z1  & \u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx64792z1 ),
	.datab(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y11_N26
cycloneii_lcell_comb \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_14_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  & \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10  & VCC # 
// !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  & 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx253z1  & (!\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1 ))

	.dataa(\u_fir|tap_array_14_filter_block_next_sum_add16_0|nx253z1 ),
	.datab(\u_fir|tap_array_15_filter_block_prod_mults28_0|nx15210z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_15_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N24
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|taps_16__15_  $ \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx64792z1  $ !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z13 ) # GND
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx64792z1  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z13 ) # !\u_fir|taps_16__15_  & 
// \u_fir|tap_array_15_filter_block_next_sum_add16_0|nx64792z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|taps_16__15_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx64792z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X45_Y14_N26
cycloneii_lcell_comb \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1  = \u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10  & VCC # 
// !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|taps_16__15_  & (\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1  & 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|taps_16__15_  & !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|taps_16__15_  & 
// (!\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1 ))

	.dataa(\u_fir|taps_16__15_ ),
	.datab(\u_fir|tap_array_15_filter_block_next_sum_add16_0|nx253z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_16_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N24
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52927 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx64792z1  = (\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z1  $ \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx64792z1  $ !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z13 ) # 
// GND
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10  = CARRY(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z1  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx64792z1  # !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z13 
// ) # !\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z1  & \u_fir|tap_array_16_filter_block_next_sum_add16_0|nx64792z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z13 )

	.dataa(\u_fir|tap_array_17_filter_block_prod_mults28_0|nx12219z1 ),
	.datab(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx64792z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z13 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx64792z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52927 .lut_mask = 16'h698E;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X42_Y14_N26
cycloneii_lcell_comb \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52926 (
// Equation(s):
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx253z1  = \u_fir|tap_array_17_filter_block_tap_next_15_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1  & \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10  & VCC # 
// !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10 ) # !\u_fir|tap_array_17_filter_block_tap_next_15_  & (\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1  & 
// !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1  & (\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10  # GND))
// \u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z7  = CARRY(\u_fir|tap_array_17_filter_block_tap_next_15_  & !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1  & !\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10  # 
// !\u_fir|tap_array_17_filter_block_tap_next_15_  & (!\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10  # !\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1 ))

	.dataa(\u_fir|tap_array_17_filter_block_tap_next_15_ ),
	.datab(\u_fir|tap_array_16_filter_block_next_sum_add16_0|nx253z1 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z10 ),
	.combout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx253z1 ),
	.cout(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx2247z7 ));
// synopsys translate_off
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52926 .lut_mask = 16'h9617;
defparam \u_fir|tap_array_17_filter_block_next_sum_add16_0|ix2247z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X35_Y14_N19
cycloneii_lcell_ff reg_audio_out_13_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\audio_out_13_~feeder_combout ),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx253z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_13_));

// atom is at LCCOMB_X35_Y14_N12
cycloneii_lcell_comb \audio_out_12_~feeder (
// Equation(s):
// \audio_out_12_~feeder_combout  = raw_audio_11_

	.dataa(vcc),
	.datab(raw_audio_11_),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\audio_out_12_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \audio_out_12_~feeder .lut_mask = 16'hCCCC;
defparam \audio_out_12_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X35_Y14_N13
cycloneii_lcell_ff reg_audio_out_12_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\audio_out_12_~feeder_combout ),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx64792z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_12_));

// atom is at LCCOMB_X35_Y14_N30
cycloneii_lcell_comb ix24999z52932(
// Equation(s):
// nx24999z9 = bit_position_0_ & (bit_position_1_ & audio_out_12_) # !bit_position_0_ & (audio_out_13_ # !bit_position_1_)

	.dataa(bit_position_0_),
	.datab(audio_out_13_),
	.datac(bit_position_1_),
	.datad(audio_out_12_),
	.cin(gnd),
	.combout(nx24999z9),
	.cout());
// synopsys translate_off
defparam ix24999z52932.lut_mask = 16'hE545;
defparam ix24999z52932.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X35_Y14_N0
cycloneii_lcell_comb \audio_out_14_~feeder (
// Equation(s):
// \audio_out_14_~feeder_combout  = raw_audio_11_

	.dataa(vcc),
	.datab(raw_audio_11_),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\audio_out_14_~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \audio_out_14_~feeder .lut_mask = 16'hCCCC;
defparam \audio_out_14_~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X35_Y14_N1
cycloneii_lcell_ff reg_audio_out_14_(
	.clk(\aud_adclrck_dup0~clkctrl_outclk ),
	.datain(\audio_out_14_~feeder_combout ),
	.sdata(\u_fir|tap_array_17_filter_block_next_sum_add16_0|nx1250z1 ),
	.aclr(gnd),
	.sclr(gnd),
	.sload(\sw~combout [16]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(audio_out_14_));

// atom is at LCCOMB_X35_Y14_N28
cycloneii_lcell_comb ix24999z52931(
// Equation(s):
// nx24999z8 = nx24999z9 & (audio_out_15_ # bit_position_1_) # !nx24999z9 & (!bit_position_1_ & audio_out_14_)

	.dataa(audio_out_15_),
	.datab(nx24999z9),
	.datac(bit_position_1_),
	.datad(audio_out_14_),
	.cin(gnd),
	.combout(nx24999z8),
	.cout());
// synopsys translate_off
defparam ix24999z52931.lut_mask = 16'hCBC8;
defparam ix24999z52931.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X35_Y14_N6
cycloneii_lcell_comb ix24999z52923(
// Equation(s):
// aud_dacdat_dup0 = bit_position_3_ & (nx24999z1) # !bit_position_3_ & (nx24999z1 & (nx24999z8) # !nx24999z1 & nx24999z6)

	.dataa(bit_position_3_),
	.datab(nx24999z6),
	.datac(nx24999z1),
	.datad(nx24999z8),
	.cin(gnd),
	.combout(aud_dacdat_dup0),
	.cout());
// synopsys translate_off
defparam ix24999z52923.lut_mask = 16'hF4A4;
defparam ix24999z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N12
cycloneii_lcell_comb \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52929 (
// Equation(s):
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx51271z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  $ VCC
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z10  = CARRY(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx51271z1 ),
	.cout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z10 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52929 .lut_mask = 16'h55AA;
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52929 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N14
cycloneii_lcell_comb \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52928 (
// Equation(s):
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx52268z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z10  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & 
// (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z10  # GND)
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z8  = CARRY(!\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z10  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z10 ),
	.combout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx52268z1 ),
	.cout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z8 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52928 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y19_N0
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52939 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx51271z1  = \u_i2c_av_config|modgen_counter_cont|q_0_  $ VCC
// \u_i2c_av_config|modgen_counter_cont|nx22081z16  = CARRY(\u_i2c_av_config|modgen_counter_cont|q_0_ )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_0_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx51271z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z16 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52939 .lut_mask = 16'h33CC;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52939 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X54_Y19_N20
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52929 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx17096z1  = \u_i2c_av_config|modgen_counter_cont|q_10_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z7  $ GND) # !\u_i2c_av_config|modgen_counter_cont|q_10_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z7  & VCC
// \u_i2c_av_config|modgen_counter_cont|nx22081z6  = CARRY(\u_i2c_av_config|modgen_counter_cont|q_10_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z7 )

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_10_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z7 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx17096z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z6 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52929 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N21
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_10_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx17096z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_10_ ));

// atom is at LCCOMB_X54_Y19_N16
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52931 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx59247z1  = \u_i2c_av_config|modgen_counter_cont|q_8_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z9  $ GND) # !\u_i2c_av_config|modgen_counter_cont|q_8_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z9  & VCC
// \u_i2c_av_config|modgen_counter_cont|nx22081z8  = CARRY(\u_i2c_av_config|modgen_counter_cont|q_8_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z9 )

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_8_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z9 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx59247z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z8 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52931 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N17
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_8_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx59247z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_8_ ));

// atom is at LCCOMB_X55_Y19_N16
cycloneii_lcell_comb \u_i2c_av_config|ix35560z52925 (
// Equation(s):
// \u_i2c_av_config|nx35560z3  = \u_i2c_av_config|modgen_counter_cont|q_11_  & \u_i2c_av_config|modgen_counter_cont|q_9_  & \u_i2c_av_config|modgen_counter_cont|q_10_  & \u_i2c_av_config|modgen_counter_cont|q_8_ 

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_11_ ),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_9_ ),
	.datac(\u_i2c_av_config|modgen_counter_cont|q_10_ ),
	.datad(\u_i2c_av_config|modgen_counter_cont|q_8_ ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx35560z3 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix35560z52925 .lut_mask = 16'h8000;
defparam \u_i2c_av_config|ix35560z52925 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X54_Y19_N6
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52936 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx54262z1  = \u_i2c_av_config|modgen_counter_cont|q_3_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z14  # !\u_i2c_av_config|modgen_counter_cont|q_3_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z14  # GND)
// \u_i2c_av_config|modgen_counter_cont|nx22081z13  = CARRY(!\u_i2c_av_config|modgen_counter_cont|nx22081z14  # !\u_i2c_av_config|modgen_counter_cont|q_3_ )

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_3_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z14 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx54262z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z13 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52936 .lut_mask = 16'h5A5F;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52936 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N7
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_3_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx54262z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_3_ ));

// atom is at LCCOMB_X55_Y19_N28
cycloneii_lcell_comb \u_i2c_av_config|ix17807z52924 (
// Equation(s):
// \u_i2c_av_config|nx17807z2  = \u_i2c_av_config|modgen_counter_cont|q_0_  & \u_i2c_av_config|modgen_counter_cont|q_3_  & \u_i2c_av_config|modgen_counter_cont|q_2_  & \u_i2c_av_config|modgen_counter_cont|q_1_ 

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_0_ ),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_3_ ),
	.datac(\u_i2c_av_config|modgen_counter_cont|q_2_ ),
	.datad(\u_i2c_av_config|modgen_counter_cont|q_1_ ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx17807z2 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix17807z52924 .lut_mask = 16'h8000;
defparam \u_i2c_av_config|ix17807z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X55_Y19_N4
cycloneii_lcell_comb \u_i2c_av_config|ix35560z52923 (
// Equation(s):
// \u_i2c_av_config|nx35560z1  = !\u_i2c_av_config|nx17807z2  # !\u_i2c_av_config|nx35560z3  # !\u_i2c_av_config|nx35560z4  # !\u_i2c_av_config|nx35560z2 

	.dataa(\u_i2c_av_config|nx35560z2 ),
	.datab(\u_i2c_av_config|nx35560z4 ),
	.datac(\u_i2c_av_config|nx35560z3 ),
	.datad(\u_i2c_av_config|nx17807z2 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx35560z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix35560z52923 .lut_mask = 16'h7FFF;
defparam \u_i2c_av_config|ix35560z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N1
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_0_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx51271z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_0_ ));

// atom is at LCCOMB_X54_Y19_N2
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52938 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx52268z1  = \u_i2c_av_config|modgen_counter_cont|q_1_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z16  # !\u_i2c_av_config|modgen_counter_cont|q_1_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z16  # GND)
// \u_i2c_av_config|modgen_counter_cont|nx22081z15  = CARRY(!\u_i2c_av_config|modgen_counter_cont|nx22081z16  # !\u_i2c_av_config|modgen_counter_cont|q_1_ )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z16 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx52268z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z15 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52938 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52938 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N3
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_1_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx52268z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_1_ ));

// atom is at LCCOMB_X54_Y19_N4
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52937 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx53265z1  = \u_i2c_av_config|modgen_counter_cont|q_2_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z15  $ GND) # !\u_i2c_av_config|modgen_counter_cont|q_2_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z15  & VCC
// \u_i2c_av_config|modgen_counter_cont|nx22081z14  = CARRY(\u_i2c_av_config|modgen_counter_cont|q_2_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z15 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_2_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z15 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx53265z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z14 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52937 .lut_mask = 16'hC30C;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52937 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N5
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_2_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx53265z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_2_ ));

// atom is at LCCOMB_X54_Y19_N8
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52935 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx55259z1  = \u_i2c_av_config|modgen_counter_cont|q_4_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z13  $ GND) # !\u_i2c_av_config|modgen_counter_cont|q_4_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z13  & VCC
// \u_i2c_av_config|modgen_counter_cont|nx22081z12  = CARRY(\u_i2c_av_config|modgen_counter_cont|q_4_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z13 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_4_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z13 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx55259z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z12 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52935 .lut_mask = 16'hC30C;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52935 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N9
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_4_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx55259z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_4_ ));

// atom is at LCCOMB_X54_Y19_N14
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52932 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx58250z1  = \u_i2c_av_config|modgen_counter_cont|q_7_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z10  # !\u_i2c_av_config|modgen_counter_cont|q_7_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z10  # GND)
// \u_i2c_av_config|modgen_counter_cont|nx22081z9  = CARRY(!\u_i2c_av_config|modgen_counter_cont|nx22081z10  # !\u_i2c_av_config|modgen_counter_cont|q_7_ )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_7_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z10 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx58250z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z9 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52932 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52932 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N15
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_7_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx58250z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_7_ ));

// atom is at LCCOMB_X54_Y19_N18
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52930 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx60244z1  = \u_i2c_av_config|modgen_counter_cont|q_9_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z8  # !\u_i2c_av_config|modgen_counter_cont|q_9_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z8  # GND)
// \u_i2c_av_config|modgen_counter_cont|nx22081z7  = CARRY(!\u_i2c_av_config|modgen_counter_cont|nx22081z8  # !\u_i2c_av_config|modgen_counter_cont|q_9_ )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_9_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z8 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx60244z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z7 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52930 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52930 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N19
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_9_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx60244z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_9_ ));

// atom is at LCCOMB_X54_Y19_N22
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52928 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx18093z1  = \u_i2c_av_config|modgen_counter_cont|q_11_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z6  # !\u_i2c_av_config|modgen_counter_cont|q_11_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z6  # GND)
// \u_i2c_av_config|modgen_counter_cont|nx22081z5  = CARRY(!\u_i2c_av_config|modgen_counter_cont|nx22081z6  # !\u_i2c_av_config|modgen_counter_cont|q_11_ )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_11_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z6 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx18093z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z5 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52928 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N23
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_11_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx18093z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_11_ ));

// atom is at LCCOMB_X54_Y19_N24
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52927 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx19090z1  = \u_i2c_av_config|modgen_counter_cont|q_12_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z5  $ GND) # !\u_i2c_av_config|modgen_counter_cont|q_12_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z5  & VCC
// \u_i2c_av_config|modgen_counter_cont|nx22081z4  = CARRY(\u_i2c_av_config|modgen_counter_cont|q_12_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z5 )

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_12_ ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z5 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx19090z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z4 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52927 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X54_Y19_N26
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52926 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx20087z1  = \u_i2c_av_config|modgen_counter_cont|q_13_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z4  # !\u_i2c_av_config|modgen_counter_cont|q_13_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z4  # GND)
// \u_i2c_av_config|modgen_counter_cont|nx22081z3  = CARRY(!\u_i2c_av_config|modgen_counter_cont|nx22081z4  # !\u_i2c_av_config|modgen_counter_cont|q_13_ )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_13_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z4 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx20087z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z3 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52926 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N27
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_13_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx20087z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_13_ ));

// atom is at LCCOMB_X54_Y19_N28
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52925 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx21084z1  = \u_i2c_av_config|modgen_counter_cont|q_14_  & (\u_i2c_av_config|modgen_counter_cont|nx22081z3  $ GND) # !\u_i2c_av_config|modgen_counter_cont|q_14_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z3  & VCC
// \u_i2c_av_config|modgen_counter_cont|nx22081z2  = CARRY(\u_i2c_av_config|modgen_counter_cont|q_14_  & !\u_i2c_av_config|modgen_counter_cont|nx22081z3 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_14_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z3 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx21084z1 ),
	.cout(\u_i2c_av_config|modgen_counter_cont|nx22081z2 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52925 .lut_mask = 16'hC30C;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N29
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_14_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx21084z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_14_ ));

// atom is at LCCOMB_X54_Y19_N30
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_cont|ix22081z52923 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_cont|nx22081z1  = \u_i2c_av_config|modgen_counter_cont|nx22081z2  $ \u_i2c_av_config|modgen_counter_cont|q_15_ 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_i2c_av_config|modgen_counter_cont|q_15_ ),
	.cin(\u_i2c_av_config|modgen_counter_cont|nx22081z2 ),
	.combout(\u_i2c_av_config|modgen_counter_cont|nx22081z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52923 .lut_mask = 16'h0FF0;
defparam \u_i2c_av_config|modgen_counter_cont|ix22081z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X54_Y19_N31
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_15_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx22081z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_15_ ));

// atom is at LCFF_X54_Y19_N25
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_cont|reg_q_12_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_cont|nx19090z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\u_i2c_av_config|nx35560z1 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_cont|q_12_ ));

// atom is at LCCOMB_X55_Y19_N2
cycloneii_lcell_comb \u_i2c_av_config|ix35560z52926 (
// Equation(s):
// \u_i2c_av_config|nx35560z4  = \u_i2c_av_config|modgen_counter_cont|q_14_  & \u_i2c_av_config|modgen_counter_cont|q_13_  & \u_i2c_av_config|modgen_counter_cont|q_15_  & \u_i2c_av_config|modgen_counter_cont|q_12_ 

	.dataa(\u_i2c_av_config|modgen_counter_cont|q_14_ ),
	.datab(\u_i2c_av_config|modgen_counter_cont|q_13_ ),
	.datac(\u_i2c_av_config|modgen_counter_cont|q_15_ ),
	.datad(\u_i2c_av_config|modgen_counter_cont|q_12_ ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx35560z4 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix35560z52926 .lut_mask = 16'h8000;
defparam \u_i2c_av_config|ix35560z52926 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X55_Y19_N18
cycloneii_lcell_comb \u_i2c_av_config|ix17807z52923 (
// Equation(s):
// \u_i2c_av_config|nx17807z1  = \u_i2c_av_config|nx35560z2  & \u_i2c_av_config|nx35560z4  & \u_i2c_av_config|nx35560z3  & \u_i2c_av_config|nx17807z2 

	.dataa(\u_i2c_av_config|nx35560z2 ),
	.datab(\u_i2c_av_config|nx35560z4 ),
	.datac(\u_i2c_av_config|nx35560z3 ),
	.datad(\u_i2c_av_config|nx17807z2 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx17807z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix17807z52923 .lut_mask = 16'h8000;
defparam \u_i2c_av_config|ix17807z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X55_Y19_N19
cycloneii_lcell_ff \u_i2c_av_config|reg_reset_n (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|nx17807z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|reset_n ));

// atom is at LCCOMB_X60_Y19_N4
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52936 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx51271z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z25  $ VCC
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z24  = CARRY(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z25 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z25 ),
	.datac(vcc),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx51271z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z24 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52936 .lut_mask = 16'h33CC;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52936 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N4
cycloneii_lcell_comb \u_i2c_av_config|ix23875z52923 (
// Equation(s):
// \u_i2c_av_config|nx23875z1  = \u_i2c_av_config|nx2692z2  # !\u_i2c_av_config|reset_n 

	.dataa(vcc),
	.datab(vcc),
	.datac(\u_i2c_av_config|reset_n ),
	.datad(\u_i2c_av_config|nx2692z2 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx23875z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix23875z52923 .lut_mask = 16'hFF0F;
defparam \u_i2c_av_config|ix23875z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N5
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_0_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx51271z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z25 ));

// atom is at LCCOMB_X60_Y19_N8
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52934 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx53265z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z21  & (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z22  $ GND) # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z21  & 
// !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z22  & VCC
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z20  = CARRY(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z21  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z22 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z21 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z22 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx53265z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z20 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52934 .lut_mask = 16'hC30C;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52934 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N9
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_2_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx53265z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z21 ));

// atom is at LCCOMB_X60_Y19_N10
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52933 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx54262z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z19  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z20  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z19  & 
// (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z20  # GND)
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z18  = CARRY(!\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z20  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z19 )

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z19 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z20 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx54262z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z18 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52933 .lut_mask = 16'h5A5F;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52933 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X60_Y19_N14
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52931 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx56256z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z15  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z16  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z15  & 
// (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z16  # GND)
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z14  = CARRY(!\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z16  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z15 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z15 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z16 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx56256z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z14 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52931 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52931 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N15
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_5_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx56256z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z15 ));

// atom is at LCCOMB_X60_Y19_N18
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52929 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx58250z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z11  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z12  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z11  & 
// (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z12  # GND)
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z10  = CARRY(!\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z12  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z11 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z11 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z12 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx58250z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z10 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52929 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52929 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N19
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_7_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx58250z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z11 ));

// atom is at LCCOMB_X60_Y19_N20
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52928 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx59247z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z9  & (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z10  $ GND) # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z9  & 
// !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z10  & VCC
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z8  = CARRY(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z9  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z10 )

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z9 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z10 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx59247z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z8 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52928 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52928 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N21
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_8_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx59247z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z9 ));

// atom is at LCCOMB_X60_Y19_N22
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52927 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx60244z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z7  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z8  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z7  & 
// (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z8  # GND)
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z6  = CARRY(!\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z8  # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z7 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z7 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z8 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx60244z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z6 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52927 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N23
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_9_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx60244z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z7 ));

// atom is at LCCOMB_X60_Y19_N24
cycloneii_lcell_comb \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52926 (
// Equation(s):
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx17096z1  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z5  & (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z6  $ GND) # !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z5  & 
// !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z6  & VCC
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z4  = CARRY(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z5  & !\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z6 )

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z5 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z6 ),
	.combout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx17096z1 ),
	.cout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z4 ));
// synopsys translate_off
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52926 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|modgen_counter_m_i2c_clk_div|ix19090z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N27
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_11_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx18093z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3 ));

// atom is at LCCOMB_X59_Y19_N26
cycloneii_lcell_comb \u_i2c_av_config|ix2692z52926 (
// Equation(s):
// \u_i2c_av_config|nx2692z4  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z13  & \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z9  & \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3  & 
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z11 

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z13 ),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z9 ),
	.datac(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3 ),
	.datad(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z11 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx2692z4 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix2692z52926 .lut_mask = 16'h8000;
defparam \u_i2c_av_config|ix2692z52926 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N11
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_3_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx54262z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z19 ));

// atom is at LCCOMB_X59_Y19_N24
cycloneii_lcell_comb \u_i2c_av_config|ix2692z52925 (
// Equation(s):
// \u_i2c_av_config|nx2692z3  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z17  # \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z19  # \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z15  # 
// \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z21 

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z17 ),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z19 ),
	.datac(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z15 ),
	.datad(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z21 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx2692z3 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix2692z52925 .lut_mask = 16'hFFFE;
defparam \u_i2c_av_config|ix2692z52925 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X60_Y19_N25
cycloneii_lcell_ff \u_i2c_av_config|modgen_counter_m_i2c_clk_div|reg_q_10_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx17096z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(\u_i2c_av_config|nx23875z1 ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z5 ));

// atom is at LCCOMB_X59_Y19_N28
cycloneii_lcell_comb \u_i2c_av_config|ix2692z52927 (
// Equation(s):
// \u_i2c_av_config|nx2692z5  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3  & (\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z7  # \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z5 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z7 ),
	.datac(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z3 ),
	.datad(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx19090z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx2692z5 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix2692z52927 .lut_mask = 16'hF0C0;
defparam \u_i2c_av_config|ix2692z52927 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N30
cycloneii_lcell_comb \u_i2c_av_config|ix2692z52924 (
// Equation(s):
// \u_i2c_av_config|nx2692z2  = \u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx1963z1  # \u_i2c_av_config|nx2692z5  # \u_i2c_av_config|nx2692z4  & \u_i2c_av_config|nx2692z3 

	.dataa(\u_i2c_av_config|modgen_counter_m_i2c_clk_div|nx1963z1 ),
	.datab(\u_i2c_av_config|nx2692z4 ),
	.datac(\u_i2c_av_config|nx2692z3 ),
	.datad(\u_i2c_av_config|nx2692z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx2692z2 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix2692z52924 .lut_mask = 16'hFFEA;
defparam \u_i2c_av_config|ix2692z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X55_Y19_N24
cycloneii_lcell_comb \u_i2c_av_config|ix2692z52923 (
// Equation(s):
// \u_i2c_av_config|nx2692z1  = \u_i2c_av_config|m_i2c_ctrl_clk  $ \u_i2c_av_config|nx2692z2 

	.dataa(vcc),
	.datab(vcc),
	.datac(\u_i2c_av_config|m_i2c_ctrl_clk ),
	.datad(\u_i2c_av_config|nx2692z2 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx2692z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix2692z52923 .lut_mask = 16'h0FF0;
defparam \u_i2c_av_config|ix2692z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X55_Y19_N25
cycloneii_lcell_ff \u_i2c_av_config|reg_m_i2c_ctrl_clk (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|nx2692z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(!\u_i2c_av_config|reset_n ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|m_i2c_ctrl_clk ));

// atom is at LCCOMB_X59_Y19_N20
cycloneii_lcell_comb \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52925 (
// Equation(s):
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  & (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z4  $ GND) # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  & 
// !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z4  & VCC
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z2  = CARRY(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z4 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z4 ),
	.combout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z1 ),
	.cout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z2 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52925 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52925 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N22
cycloneii_lcell_comb \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52923 (
// Equation(s):
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z2  $ \u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.cin(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z2 ),
	.combout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52923 .lut_mask = 16'h0FF0;
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X59_Y19_N23
cycloneii_lcell_ff \u_i2c_av_config|u0|modgen_counter_sd_counter|reg_q_5_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z1 ),
	.sdata(vcc),
	.aclr(gnd),
	.sclr(gnd),
	.sload(!\u_i2c_av_config|reset_n ),
	.ena(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ));

// atom is at LCFF_X59_Y19_N13
cycloneii_lcell_ff \u_i2c_av_config|u0|modgen_counter_sd_counter|reg_q_0_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx51271z1 ),
	.sdata(vcc),
	.aclr(gnd),
	.sclr(gnd),
	.sload(!\u_i2c_av_config|reset_n ),
	.ena(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ));

// atom is at LCCOMB_X59_Y19_N8
cycloneii_lcell_comb \u_i2c_av_config|u0|ix7286z52923 (
// Equation(s):
// \u_i2c_av_config|u0|nx7286z1  = \u_i2c_av_config|u0|nx7286z2  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 

	.dataa(\u_i2c_av_config|u0|nx7286z2 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datac(vcc),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx7286z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix7286z52923 .lut_mask = 16'hBBFF;
defparam \u_i2c_av_config|u0|ix7286z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N0
cycloneii_lcell_comb \u_i2c_av_config|ix51161z52923 (
// Equation(s):
// \u_i2c_av_config|nx51161z1  = \u_i2c_av_config|reset_n  & (\u_i2c_av_config|m_i2c_ctrl_clk  $ \u_i2c_av_config|nx2692z2 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|m_i2c_ctrl_clk ),
	.datac(\u_i2c_av_config|reset_n ),
	.datad(\u_i2c_av_config|nx2692z2 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|nx51161z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|ix51161z52923 .lut_mask = 16'h30C0;
defparam \u_i2c_av_config|ix51161z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N2
cycloneii_lcell_comb \u_i2c_av_config|u0|modgen_counter_sd_counter|ix55259z52924 (
// Equation(s):
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3  = !\u_i2c_av_config|m_i2c_ctrl_clk  & \u_i2c_av_config|nx51161z1  & (\u_i2c_av_config|u0|nx7286z1  # !\u_i2c_av_config|reset_n )

	.dataa(\u_i2c_av_config|reset_n ),
	.datab(\u_i2c_av_config|m_i2c_ctrl_clk ),
	.datac(\u_i2c_av_config|u0|nx7286z1 ),
	.datad(\u_i2c_av_config|nx51161z1 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix55259z52924 .lut_mask = 16'h3100;
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix55259z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X59_Y19_N15
cycloneii_lcell_ff \u_i2c_av_config|u0|modgen_counter_sd_counter|reg_q_1_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx52268z1 ),
	.sdata(vcc),
	.aclr(gnd),
	.sclr(gnd),
	.sload(!\u_i2c_av_config|reset_n ),
	.ena(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ));

// atom is at LCCOMB_X59_Y19_N16
cycloneii_lcell_comb \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52927 (
// Equation(s):
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx53265z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z8  $ GND) # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & 
// !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z8  & VCC
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z6  = CARRY(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z8 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datab(vcc),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z8 ),
	.combout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx53265z1 ),
	.cout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z6 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52927 .lut_mask = 16'hA50A;
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N18
cycloneii_lcell_comb \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52926 (
// Equation(s):
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx54262z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z6  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  & 
// (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z6  # GND)
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z4  = CARRY(!\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z6  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 )

	.dataa(vcc),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z6 ),
	.combout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx54262z1 ),
	.cout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z4 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52926 .lut_mask = 16'h3C3F;
defparam \u_i2c_av_config|u0|modgen_counter_sd_counter|ix56256z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCFF_X59_Y19_N19
cycloneii_lcell_ff \u_i2c_av_config|u0|modgen_counter_sd_counter|reg_q_3_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx54262z1 ),
	.sdata(vcc),
	.aclr(gnd),
	.sclr(gnd),
	.sload(!\u_i2c_av_config|reset_n ),
	.ena(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ));

// atom is at LCFF_X59_Y19_N21
cycloneii_lcell_ff \u_i2c_av_config|u0|modgen_counter_sd_counter|reg_q_4_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z1 ),
	.sdata(vcc),
	.aclr(gnd),
	.sclr(gnd),
	.sload(!\u_i2c_av_config|reset_n ),
	.ena(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ));

// atom is at LCFF_X59_Y19_N17
cycloneii_lcell_ff \u_i2c_av_config|u0|modgen_counter_sd_counter|reg_q_2_ (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx53265z1 ),
	.sdata(vcc),
	.aclr(gnd),
	.sclr(gnd),
	.sload(!\u_i2c_av_config|reset_n ),
	.ena(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx55259z3 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ));

// atom is at LCCOMB_X57_Y19_N24
cycloneii_lcell_comb \u_i2c_av_config|u0|ix43379z52924 (
// Equation(s):
// \u_i2c_av_config|u0|nx43379z2  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  # 
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx43379z2 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix43379z52924 .lut_mask = 16'h0504;
defparam \u_i2c_av_config|u0|ix43379z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y19_N2
cycloneii_lcell_comb \u_i2c_av_config|u0|ix43379z52926 (
// Equation(s):
// \u_i2c_av_config|u0|nx43379z4  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx43379z4 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix43379z52926 .lut_mask = 16'h8080;
defparam \u_i2c_av_config|u0|ix43379z52926 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y19_N28
cycloneii_lcell_comb \u_i2c_av_config|u0|ix43379z52925 (
// Equation(s):
// \u_i2c_av_config|u0|nx43379z3  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  & (!\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  # !\u_i2c_av_config|u0|nx43379z4 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datab(\u_i2c_av_config|u0|nx43379z4 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx43379z3 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix43379z52925 .lut_mask = 16'h020A;
defparam \u_i2c_av_config|u0|ix43379z52925 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N24
cycloneii_lcell_comb \u_i2c_av_config|u0|ix44942z52923 (
// Equation(s):
// \u_i2c_av_config|u0|nx44942z1  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 

	.dataa(vcc),
	.datab(vcc),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx44942z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix44942z52923 .lut_mask = 16'h0F00;
defparam \u_i2c_av_config|u0|ix44942z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N18
cycloneii_lcell_comb \u_i2c_av_config|u0|ix44942z52929 (
// Equation(s):
// \u_i2c_av_config|u0|nx44942z7  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx44942z7 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix44942z52929 .lut_mask = 16'h55FF;
defparam \u_i2c_av_config|u0|ix44942z52929 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N4
cycloneii_lcell_comb \u_i2c_av_config|u0|ix44942z52928 (
// Equation(s):
// \u_i2c_av_config|u0|nx44942z6  = !\u_i2c_av_config|u0|nx44942z8  & !\u_i2c_av_config|u0|nx44942z7  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  # !\u_i2c_av_config|reset_n 

	.dataa(\u_i2c_av_config|u0|nx44942z8 ),
	.datab(\u_i2c_av_config|u0|nx44942z7 ),
	.datac(\u_i2c_av_config|reset_n ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx44942z6 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix44942z52928 .lut_mask = 16'h0F1F;
defparam \u_i2c_av_config|u0|ix44942z52928 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N26
cycloneii_lcell_comb \u_i2c_av_config|u0|ix44942z52927 (
// Equation(s):
// \u_i2c_av_config|u0|nx44942z5  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  # \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 

	.dataa(vcc),
	.datab(vcc),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx44942z5 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix44942z52927 .lut_mask = 16'hFFF0;
defparam \u_i2c_av_config|u0|ix44942z52927 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N14
cycloneii_lcell_comb \u_i2c_av_config|u0|ix44942z52925 (
// Equation(s):
// \u_i2c_av_config|u0|nx44942z3  = \u_i2c_av_config|u0|nx44942z6  # !\u_i2c_av_config|u0|nx44942z4  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11  & !\u_i2c_av_config|u0|nx44942z5 

	.dataa(\u_i2c_av_config|u0|nx44942z4 ),
	.datab(\u_i2c_av_config|u0|nx44942z6 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z11 ),
	.datad(\u_i2c_av_config|u0|nx44942z5 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx44942z3 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix44942z52925 .lut_mask = 16'hCCCD;
defparam \u_i2c_av_config|u0|ix44942z52925 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N8
cycloneii_lcell_comb \u_i2c_av_config|u0|ix44942z52924 (
// Equation(s):
// \u_i2c_av_config|u0|nx44942z2  = \u_i2c_av_config|u0|nx44942z3  & \u_i2c_av_config|nx51161z1  & !\u_i2c_av_config|m_i2c_ctrl_clk 

	.dataa(vcc),
	.datab(\u_i2c_av_config|u0|nx44942z3 ),
	.datac(\u_i2c_av_config|nx51161z1 ),
	.datad(\u_i2c_av_config|m_i2c_ctrl_clk ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx44942z2 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix44942z52924 .lut_mask = 16'h00C0;
defparam \u_i2c_av_config|u0|ix44942z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X58_Y19_N25
cycloneii_lcell_ff \u_i2c_av_config|u0|reg_sclk (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|u0|nx44942z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(!\u_i2c_av_config|reset_n ),
	.sload(gnd),
	.ena(\u_i2c_av_config|u0|nx44942z2 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|u0|nx43379z1 ));

// atom is at LCCOMB_X57_Y19_N6
cycloneii_lcell_comb \u_i2c_av_config|u0|ix43379z52923 (
// Equation(s):
// \u_i2c_av_config|u0|p_i2c_sclk  = !\u_i2c_av_config|m_i2c_ctrl_clk  & (\u_i2c_av_config|u0|nx43379z2  # \u_i2c_av_config|u0|nx43379z3 ) # !\u_i2c_av_config|u0|nx43379z1 

	.dataa(\u_i2c_av_config|u0|nx43379z2 ),
	.datab(\u_i2c_av_config|u0|nx43379z3 ),
	.datac(\u_i2c_av_config|m_i2c_ctrl_clk ),
	.datad(\u_i2c_av_config|u0|nx43379z1 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|p_i2c_sclk ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix43379z52923 .lut_mask = 16'h0EFF;
defparam \u_i2c_av_config|u0|ix43379z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at CLKCTRL_G9
cycloneii_clkctrl \clock_27~clkctrl (
	.ena(vcc),
	.inclk({gnd,gnd,gnd,\clock_27~combout }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\clock_27~clkctrl_outclk ));
// synopsys translate_off
defparam \clock_27~clkctrl .clock_type = "global clock";
defparam \clock_27~clkctrl .ena_register_mode = "falling edge";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N14
cycloneii_lcell_comb \u_i2c_av_config|u0|ix22137z52924 (
// Equation(s):
// \u_i2c_av_config|u0|sdo_5n5s2f1_1_  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  & (!\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  # 
// !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|sdo_5n5s2f1_1_ ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix22137z52924 .lut_mask = 16'h1115;
defparam \u_i2c_av_config|u0|ix22137z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N2
cycloneii_lcell_comb \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52927 (
// Equation(s):
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & (\u_i2c_av_config|u0|sdo_5n5s2f1_1_  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11  # !\u_i2c_av_config|u0|sdo_5n5s2f1_1_  & 
// (\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11  # GND)) # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & (\u_i2c_av_config|u0|sdo_5n5s2f1_1_  & \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11  & VCC # !\u_i2c_av_config|u0|sdo_5n5s2f1_1_  & 
// !\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11 )
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z8  = CARRY(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & (!\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11  # !\u_i2c_av_config|u0|sdo_5n5s2f1_1_ ) # 
// !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  & !\u_i2c_av_config|u0|sdo_5n5s2f1_1_  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datab(\u_i2c_av_config|u0|sdo_5n5s2f1_1_ ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z11 ),
	.combout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1 ),
	.cout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z8 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52927 .lut_mask = 16'h692B;
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52927 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N4
cycloneii_lcell_comb \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52926 (
// Equation(s):
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1  = (\u_i2c_av_config|u0|nx22137z1  $ \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  $ \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z8 ) # GND
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z5  = CARRY(\u_i2c_av_config|u0|nx22137z1  & (!\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z8  # !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ) # !\u_i2c_av_config|u0|nx22137z1  & 
// !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z8 )

	.dataa(\u_i2c_av_config|u0|nx22137z1 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datac(vcc),
	.datad(vcc),
	.cin(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z8 ),
	.combout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1 ),
	.cout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z5 ));
// synopsys translate_off
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52926 .lut_mask = 16'h962B;
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52926 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N8
cycloneii_lcell_comb \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52923 (
// Equation(s):
// \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1  = \u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z3  $ !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 

	.dataa(vcc),
	.datab(vcc),
	.datac(vcc),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.cin(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z3 ),
	.combout(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52923 .lut_mask = 16'hF00F;
defparam \u_i2c_av_config|u0|sdo_sub5_5i2|ix41961z52923 .sum_lutc_input = "cin";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N30
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52940 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z18  = \u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1 

	.dataa(\u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1 ),
	.datab(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1 ),
	.datac(\u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1 ),
	.datad(\u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z18 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52940 .lut_mask = 16'h0002;
defparam \u_i2c_av_config|u0|ix41315z52940 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N22
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52931 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z9  = \u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1  & !\u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1  & (\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1  # !\u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1 )

	.dataa(\u_i2c_av_config|u0|sdo_sub5_5i2|nx37973z1 ),
	.datab(\u_i2c_av_config|u0|sdo_sub5_5i2|nx41961z1 ),
	.datac(\u_i2c_av_config|u0|sdo_sub5_5i2|nx39967z1 ),
	.datad(\u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z9 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52931 .lut_mask = 16'h00D0;
defparam \u_i2c_av_config|u0|ix41315z52931 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y19_N0
cycloneii_lcell_comb \u_i2c_av_config|u0|ix44942z52926 (
// Equation(s):
// \u_i2c_av_config|u0|nx44942z4  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  # \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 

	.dataa(vcc),
	.datab(vcc),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx44942z4 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix44942z52926 .lut_mask = 16'hFFF0;
defparam \u_i2c_av_config|u0|ix44942z52926 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y19_N22
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52927 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z5  = \u_i2c_av_config|u0|nx44942z4  # \u_i2c_av_config|u0|nx43379z4  # \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7  & \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datab(\u_i2c_av_config|u0|nx44942z4 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.datad(\u_i2c_av_config|u0|nx43379z4 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z5 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52927 .lut_mask = 16'hFFEC;
defparam \u_i2c_av_config|u0|ix41315z52927 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y19_N16
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52928 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z6  = !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  & !\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  & (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9  # \u_i2c_av_config|u0|nx44942z5 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z9 ),
	.datab(\u_i2c_av_config|u0|nx44942z5 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z6 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52928 .lut_mask = 16'h000E;
defparam \u_i2c_av_config|u0|ix41315z52928 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X59_Y19_N6
cycloneii_lcell_comb \u_i2c_av_config|u0|ix22137z52923 (
// Equation(s):
// \u_i2c_av_config|u0|nx22137z1  = \u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1  # \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3  & (\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5  # 
// \u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 )

	.dataa(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z3 ),
	.datab(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z5 ),
	.datac(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx56256z7 ),
	.datad(\u_i2c_av_config|u0|modgen_counter_sd_counter|nx64583z1 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx22137z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix22137z52923 .lut_mask = 16'hFFA8;
defparam \u_i2c_av_config|u0|ix22137z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X57_Y19_N10
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52925 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z3  = \u_i2c_av_config|u0|nx41315z6  # \u_i2c_av_config|u0|nx22137z1  & !\u_i2c_av_config|u0|nx41315z4  # !\u_i2c_av_config|u0|nx22137z1  & (\u_i2c_av_config|u0|nx41315z5 )

	.dataa(\u_i2c_av_config|u0|nx41315z4 ),
	.datab(\u_i2c_av_config|u0|nx41315z5 ),
	.datac(\u_i2c_av_config|u0|nx41315z6 ),
	.datad(\u_i2c_av_config|u0|nx22137z1 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z3 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52925 .lut_mask = 16'hF5FC;
defparam \u_i2c_av_config|u0|ix41315z52925 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N16
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52930 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z8  = !\u_i2c_av_config|u0|sdo_sub5_5i2|nx40964z1  & \u_i2c_av_config|u0|nx41315z9  & \u_i2c_av_config|u0|nx41315z3 

	.dataa(\u_i2c_av_config|u0|sdo_sub5_5i2|nx40964z1 ),
	.datab(\u_i2c_av_config|u0|nx41315z9 ),
	.datac(\u_i2c_av_config|u0|nx41315z3 ),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z8 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52930 .lut_mask = 16'h4040;
defparam \u_i2c_av_config|u0|ix41315z52930 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N28
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52924 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z2  = !\u_i2c_av_config|u0|sdo_sub5_5i2|nx40964z1  & \u_i2c_av_config|u0|nx41315z3 

	.dataa(\u_i2c_av_config|u0|sdo_sub5_5i2|nx40964z1 ),
	.datab(vcc),
	.datac(\u_i2c_av_config|u0|nx41315z3 ),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z2 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52924 .lut_mask = 16'h5050;
defparam \u_i2c_av_config|u0|ix41315z52924 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N20
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52929 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z7  = \u_i2c_av_config|u0|nx41315z8  # \u_i2c_av_config|u0|nx41315z10  & \u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1  & \u_i2c_av_config|u0|nx41315z2 

	.dataa(\u_i2c_av_config|u0|nx41315z10 ),
	.datab(\u_i2c_av_config|u0|sdo_sub5_5i2|nx38970z1 ),
	.datac(\u_i2c_av_config|u0|nx41315z8 ),
	.datad(\u_i2c_av_config|u0|nx41315z2 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z7 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52929 .lut_mask = 16'hF8F0;
defparam \u_i2c_av_config|u0|ix41315z52929 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X56_Y19_N12
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52923 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z1  = !\u_i2c_av_config|u0|nx41315z11  & !\u_i2c_av_config|u0|nx41315z7  & (!\u_i2c_av_config|u0|nx41315z2  # !\u_i2c_av_config|u0|nx41315z18 )

	.dataa(\u_i2c_av_config|u0|nx41315z11 ),
	.datab(\u_i2c_av_config|u0|nx41315z18 ),
	.datac(\u_i2c_av_config|u0|nx41315z7 ),
	.datad(\u_i2c_av_config|u0|nx41315z2 ),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z1 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52923 .lut_mask = 16'h0105;
defparam \u_i2c_av_config|u0|ix41315z52923 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X58_Y19_N30
cycloneii_lcell_comb \u_i2c_av_config|u0|ix41315z52941 (
// Equation(s):
// \u_i2c_av_config|u0|nx41315z19  = \u_i2c_av_config|u0|nx41315z20  & !\u_i2c_av_config|m_i2c_ctrl_clk  & \u_i2c_av_config|nx51161z1 

	.dataa(\u_i2c_av_config|u0|nx41315z20 ),
	.datab(\u_i2c_av_config|m_i2c_ctrl_clk ),
	.datac(\u_i2c_av_config|nx51161z1 ),
	.datad(vcc),
	.cin(gnd),
	.combout(\u_i2c_av_config|u0|nx41315z19 ),
	.cout());
// synopsys translate_off
defparam \u_i2c_av_config|u0|ix41315z52941 .lut_mask = 16'h2020;
defparam \u_i2c_av_config|u0|ix41315z52941 .sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X56_Y19_N13
cycloneii_lcell_ff \u_i2c_av_config|u0|reg_sdo (
	.clk(\clock_27~clkctrl_outclk ),
	.datain(\u_i2c_av_config|u0|nx41315z1 ),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(!\u_i2c_av_config|reset_n ),
	.sload(gnd),
	.ena(\u_i2c_av_config|u0|nx41315z19 ),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(\u_i2c_av_config|u0|nx51857z1 ));

// atom is at LCCOMB_X35_Y2_N24
cycloneii_lcell_comb ix30102z52923(
// Equation(s):
// nx30102z1 = !u_audio_dac_bck_div_2_ & \key~combout [0]

	.dataa(vcc),
	.datab(vcc),
	.datac(u_audio_dac_bck_div_2_),
	.datad(\key~combout [0]),
	.cin(gnd),
	.combout(nx30102z1),
	.cout());
// synopsys translate_off
defparam ix30102z52923.lut_mask = 16'h0F00;
defparam ix30102z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X34_Y2_N14
cycloneii_lcell_comb ix30102z52924(
// Equation(s):
// nx30102z2 = u_audio_dac_bck_div_1_ & (u_audio_dac_bck_div_0_ # u_audio_dac_bck_div_2_) # !u_audio_dac_bck_div_1_ & u_audio_dac_bck_div_0_ & u_audio_dac_bck_div_2_ # !\key~combout [0]

	.dataa(\key~combout [0]),
	.datab(u_audio_dac_bck_div_1_),
	.datac(u_audio_dac_bck_div_0_),
	.datad(u_audio_dac_bck_div_2_),
	.cin(gnd),
	.combout(nx30102z2),
	.cout());
// synopsys translate_off
defparam ix30102z52924.lut_mask = 16'hFDD5;
defparam ix30102z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X35_Y2_N25
cycloneii_lcell_ff u_audio_dac_modgen_counter_bck_div_reg_q_2_(
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(nx30102z1),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nx30102z2),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_audio_dac_bck_div_2_));

// atom is at LCCOMB_X34_Y2_N0
cycloneii_lcell_comb ix32096z52923(
// Equation(s):
// nx32096z1 = \key~combout [0] & !u_audio_dac_bck_div_0_ & (!u_audio_dac_bck_div_2_ # !u_audio_dac_bck_div_1_)

	.dataa(\key~combout [0]),
	.datab(u_audio_dac_bck_div_1_),
	.datac(u_audio_dac_bck_div_0_),
	.datad(u_audio_dac_bck_div_2_),
	.cin(gnd),
	.combout(nx32096z1),
	.cout());
// synopsys translate_off
defparam ix32096z52923.lut_mask = 16'h020A;
defparam ix32096z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y2_N1
cycloneii_lcell_ff u_audio_dac_modgen_counter_bck_div_reg_q_0_(
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(nx32096z1),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_audio_dac_bck_div_0_));

// atom is at LCCOMB_X34_Y2_N26
cycloneii_lcell_comb ix31099z52923(
// Equation(s):
// nx31099z1 = \key~combout [0] & !u_audio_dac_bck_div_1_ & (!u_audio_dac_bck_div_2_ # !u_audio_dac_bck_div_0_)

	.dataa(\key~combout [0]),
	.datab(u_audio_dac_bck_div_0_),
	.datac(u_audio_dac_bck_div_1_),
	.datad(u_audio_dac_bck_div_2_),
	.cin(gnd),
	.combout(nx31099z1),
	.cout());
// synopsys translate_off
defparam ix31099z52923.lut_mask = 16'h020A;
defparam ix31099z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCCOMB_X34_Y2_N8
cycloneii_lcell_comb ix31099z52924(
// Equation(s):
// nx31099z2 = u_audio_dac_bck_div_0_ # u_audio_dac_bck_div_1_ & u_audio_dac_bck_div_2_ # !\key~combout [0]

	.dataa(\key~combout [0]),
	.datab(u_audio_dac_bck_div_1_),
	.datac(u_audio_dac_bck_div_0_),
	.datad(u_audio_dac_bck_div_2_),
	.cin(gnd),
	.combout(nx31099z2),
	.cout());
// synopsys translate_off
defparam ix31099z52924.lut_mask = 16'hFDF5;
defparam ix31099z52924.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y2_N27
cycloneii_lcell_ff u_audio_dac_modgen_counter_bck_div_reg_q_1_(
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(nx31099z1),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nx31099z2),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(u_audio_dac_bck_div_1_));

// atom is at LCCOMB_X34_Y2_N16
cycloneii_lcell_comb ix15494z52923(
// Equation(s):
// nx15494z1 = aud_bclk_dup0 $ (u_audio_dac_bck_div_2_ & (u_audio_dac_bck_div_0_ # u_audio_dac_bck_div_1_))

	.dataa(u_audio_dac_bck_div_0_),
	.datab(u_audio_dac_bck_div_1_),
	.datac(aud_bclk_dup0),
	.datad(u_audio_dac_bck_div_2_),
	.cin(gnd),
	.combout(nx15494z1),
	.cout());
// synopsys translate_off
defparam ix15494z52923.lut_mask = 16'h1EF0;
defparam ix15494z52923.sum_lutc_input = "datac";
// synopsys translate_on

// atom is at LCFF_X34_Y2_N17
cycloneii_lcell_ff u_audio_dac_reg_aud_bck(
	.clk(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.datain(nx15494z1),
	.sdata(gnd),
	.aclr(gnd),
	.sclr(!\key~combout [0]),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.regout(aud_bclk_dup0));

// atom is at PIN_AE22
cycloneii_io ledg_triBus1_0_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[0]));
// synopsys translate_off
defparam ledg_triBus1_0_.input_async_reset = "none";
defparam ledg_triBus1_0_.input_power_up = "low";
defparam ledg_triBus1_0_.input_register_mode = "none";
defparam ledg_triBus1_0_.input_sync_reset = "none";
defparam ledg_triBus1_0_.oe_async_reset = "none";
defparam ledg_triBus1_0_.oe_power_up = "low";
defparam ledg_triBus1_0_.oe_register_mode = "none";
defparam ledg_triBus1_0_.oe_sync_reset = "none";
defparam ledg_triBus1_0_.operation_mode = "output";
defparam ledg_triBus1_0_.output_async_reset = "none";
defparam ledg_triBus1_0_.output_power_up = "low";
defparam ledg_triBus1_0_.output_register_mode = "none";
defparam ledg_triBus1_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AF22
cycloneii_io ledg_triBus1_1_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[1]));
// synopsys translate_off
defparam ledg_triBus1_1_.input_async_reset = "none";
defparam ledg_triBus1_1_.input_power_up = "low";
defparam ledg_triBus1_1_.input_register_mode = "none";
defparam ledg_triBus1_1_.input_sync_reset = "none";
defparam ledg_triBus1_1_.oe_async_reset = "none";
defparam ledg_triBus1_1_.oe_power_up = "low";
defparam ledg_triBus1_1_.oe_register_mode = "none";
defparam ledg_triBus1_1_.oe_sync_reset = "none";
defparam ledg_triBus1_1_.operation_mode = "output";
defparam ledg_triBus1_1_.output_async_reset = "none";
defparam ledg_triBus1_1_.output_power_up = "low";
defparam ledg_triBus1_1_.output_register_mode = "none";
defparam ledg_triBus1_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_W19
cycloneii_io ledg_triBus1_2_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[2]));
// synopsys translate_off
defparam ledg_triBus1_2_.input_async_reset = "none";
defparam ledg_triBus1_2_.input_power_up = "low";
defparam ledg_triBus1_2_.input_register_mode = "none";
defparam ledg_triBus1_2_.input_sync_reset = "none";
defparam ledg_triBus1_2_.oe_async_reset = "none";
defparam ledg_triBus1_2_.oe_power_up = "low";
defparam ledg_triBus1_2_.oe_register_mode = "none";
defparam ledg_triBus1_2_.oe_sync_reset = "none";
defparam ledg_triBus1_2_.operation_mode = "output";
defparam ledg_triBus1_2_.output_async_reset = "none";
defparam ledg_triBus1_2_.output_power_up = "low";
defparam ledg_triBus1_2_.output_register_mode = "none";
defparam ledg_triBus1_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_V18
cycloneii_io ledg_triBus1_3_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[3]));
// synopsys translate_off
defparam ledg_triBus1_3_.input_async_reset = "none";
defparam ledg_triBus1_3_.input_power_up = "low";
defparam ledg_triBus1_3_.input_register_mode = "none";
defparam ledg_triBus1_3_.input_sync_reset = "none";
defparam ledg_triBus1_3_.oe_async_reset = "none";
defparam ledg_triBus1_3_.oe_power_up = "low";
defparam ledg_triBus1_3_.oe_register_mode = "none";
defparam ledg_triBus1_3_.oe_sync_reset = "none";
defparam ledg_triBus1_3_.operation_mode = "output";
defparam ledg_triBus1_3_.output_async_reset = "none";
defparam ledg_triBus1_3_.output_power_up = "low";
defparam ledg_triBus1_3_.output_register_mode = "none";
defparam ledg_triBus1_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_U18
cycloneii_io ledg_triBus1_4_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[4]));
// synopsys translate_off
defparam ledg_triBus1_4_.input_async_reset = "none";
defparam ledg_triBus1_4_.input_power_up = "low";
defparam ledg_triBus1_4_.input_register_mode = "none";
defparam ledg_triBus1_4_.input_sync_reset = "none";
defparam ledg_triBus1_4_.oe_async_reset = "none";
defparam ledg_triBus1_4_.oe_power_up = "low";
defparam ledg_triBus1_4_.oe_register_mode = "none";
defparam ledg_triBus1_4_.oe_sync_reset = "none";
defparam ledg_triBus1_4_.operation_mode = "output";
defparam ledg_triBus1_4_.output_async_reset = "none";
defparam ledg_triBus1_4_.output_power_up = "low";
defparam ledg_triBus1_4_.output_register_mode = "none";
defparam ledg_triBus1_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_U17
cycloneii_io ledg_triBus1_5_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[5]));
// synopsys translate_off
defparam ledg_triBus1_5_.input_async_reset = "none";
defparam ledg_triBus1_5_.input_power_up = "low";
defparam ledg_triBus1_5_.input_register_mode = "none";
defparam ledg_triBus1_5_.input_sync_reset = "none";
defparam ledg_triBus1_5_.oe_async_reset = "none";
defparam ledg_triBus1_5_.oe_power_up = "low";
defparam ledg_triBus1_5_.oe_register_mode = "none";
defparam ledg_triBus1_5_.oe_sync_reset = "none";
defparam ledg_triBus1_5_.operation_mode = "output";
defparam ledg_triBus1_5_.output_async_reset = "none";
defparam ledg_triBus1_5_.output_power_up = "low";
defparam ledg_triBus1_5_.output_register_mode = "none";
defparam ledg_triBus1_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AA20
cycloneii_io ledg_triBus1_6_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[6]));
// synopsys translate_off
defparam ledg_triBus1_6_.input_async_reset = "none";
defparam ledg_triBus1_6_.input_power_up = "low";
defparam ledg_triBus1_6_.input_register_mode = "none";
defparam ledg_triBus1_6_.input_sync_reset = "none";
defparam ledg_triBus1_6_.oe_async_reset = "none";
defparam ledg_triBus1_6_.oe_power_up = "low";
defparam ledg_triBus1_6_.oe_register_mode = "none";
defparam ledg_triBus1_6_.oe_sync_reset = "none";
defparam ledg_triBus1_6_.operation_mode = "output";
defparam ledg_triBus1_6_.output_async_reset = "none";
defparam ledg_triBus1_6_.output_power_up = "low";
defparam ledg_triBus1_6_.output_register_mode = "none";
defparam ledg_triBus1_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_Y18
cycloneii_io ledg_triBus1_7_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[7]));
// synopsys translate_off
defparam ledg_triBus1_7_.input_async_reset = "none";
defparam ledg_triBus1_7_.input_power_up = "low";
defparam ledg_triBus1_7_.input_register_mode = "none";
defparam ledg_triBus1_7_.input_sync_reset = "none";
defparam ledg_triBus1_7_.oe_async_reset = "none";
defparam ledg_triBus1_7_.oe_power_up = "low";
defparam ledg_triBus1_7_.oe_register_mode = "none";
defparam ledg_triBus1_7_.oe_sync_reset = "none";
defparam ledg_triBus1_7_.operation_mode = "output";
defparam ledg_triBus1_7_.output_async_reset = "none";
defparam ledg_triBus1_7_.output_power_up = "low";
defparam ledg_triBus1_7_.output_register_mode = "none";
defparam ledg_triBus1_7_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_Y12
cycloneii_io ledg_triBus1_8_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledg[8]));
// synopsys translate_off
defparam ledg_triBus1_8_.input_async_reset = "none";
defparam ledg_triBus1_8_.input_power_up = "low";
defparam ledg_triBus1_8_.input_register_mode = "none";
defparam ledg_triBus1_8_.input_sync_reset = "none";
defparam ledg_triBus1_8_.oe_async_reset = "none";
defparam ledg_triBus1_8_.oe_power_up = "low";
defparam ledg_triBus1_8_.oe_register_mode = "none";
defparam ledg_triBus1_8_.oe_sync_reset = "none";
defparam ledg_triBus1_8_.operation_mode = "output";
defparam ledg_triBus1_8_.output_async_reset = "none";
defparam ledg_triBus1_8_.output_power_up = "low";
defparam ledg_triBus1_8_.output_register_mode = "none";
defparam ledg_triBus1_8_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AE23
cycloneii_io ledr_triBus2_0_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[0]));
// synopsys translate_off
defparam ledr_triBus2_0_.input_async_reset = "none";
defparam ledr_triBus2_0_.input_power_up = "low";
defparam ledr_triBus2_0_.input_register_mode = "none";
defparam ledr_triBus2_0_.input_sync_reset = "none";
defparam ledr_triBus2_0_.oe_async_reset = "none";
defparam ledr_triBus2_0_.oe_power_up = "low";
defparam ledr_triBus2_0_.oe_register_mode = "none";
defparam ledr_triBus2_0_.oe_sync_reset = "none";
defparam ledr_triBus2_0_.operation_mode = "output";
defparam ledr_triBus2_0_.output_async_reset = "none";
defparam ledr_triBus2_0_.output_power_up = "low";
defparam ledr_triBus2_0_.output_register_mode = "none";
defparam ledr_triBus2_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AF23
cycloneii_io ledr_triBus2_1_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[1]));
// synopsys translate_off
defparam ledr_triBus2_1_.input_async_reset = "none";
defparam ledr_triBus2_1_.input_power_up = "low";
defparam ledr_triBus2_1_.input_register_mode = "none";
defparam ledr_triBus2_1_.input_sync_reset = "none";
defparam ledr_triBus2_1_.oe_async_reset = "none";
defparam ledr_triBus2_1_.oe_power_up = "low";
defparam ledr_triBus2_1_.oe_register_mode = "none";
defparam ledr_triBus2_1_.oe_sync_reset = "none";
defparam ledr_triBus2_1_.operation_mode = "output";
defparam ledr_triBus2_1_.output_async_reset = "none";
defparam ledr_triBus2_1_.output_power_up = "low";
defparam ledr_triBus2_1_.output_register_mode = "none";
defparam ledr_triBus2_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AB21
cycloneii_io ledr_triBus2_2_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[2]));
// synopsys translate_off
defparam ledr_triBus2_2_.input_async_reset = "none";
defparam ledr_triBus2_2_.input_power_up = "low";
defparam ledr_triBus2_2_.input_register_mode = "none";
defparam ledr_triBus2_2_.input_sync_reset = "none";
defparam ledr_triBus2_2_.oe_async_reset = "none";
defparam ledr_triBus2_2_.oe_power_up = "low";
defparam ledr_triBus2_2_.oe_register_mode = "none";
defparam ledr_triBus2_2_.oe_sync_reset = "none";
defparam ledr_triBus2_2_.operation_mode = "output";
defparam ledr_triBus2_2_.output_async_reset = "none";
defparam ledr_triBus2_2_.output_power_up = "low";
defparam ledr_triBus2_2_.output_register_mode = "none";
defparam ledr_triBus2_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AC22
cycloneii_io ledr_triBus2_3_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[3]));
// synopsys translate_off
defparam ledr_triBus2_3_.input_async_reset = "none";
defparam ledr_triBus2_3_.input_power_up = "low";
defparam ledr_triBus2_3_.input_register_mode = "none";
defparam ledr_triBus2_3_.input_sync_reset = "none";
defparam ledr_triBus2_3_.oe_async_reset = "none";
defparam ledr_triBus2_3_.oe_power_up = "low";
defparam ledr_triBus2_3_.oe_register_mode = "none";
defparam ledr_triBus2_3_.oe_sync_reset = "none";
defparam ledr_triBus2_3_.operation_mode = "output";
defparam ledr_triBus2_3_.output_async_reset = "none";
defparam ledr_triBus2_3_.output_power_up = "low";
defparam ledr_triBus2_3_.output_register_mode = "none";
defparam ledr_triBus2_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AD22
cycloneii_io ledr_triBus2_4_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[4]));
// synopsys translate_off
defparam ledr_triBus2_4_.input_async_reset = "none";
defparam ledr_triBus2_4_.input_power_up = "low";
defparam ledr_triBus2_4_.input_register_mode = "none";
defparam ledr_triBus2_4_.input_sync_reset = "none";
defparam ledr_triBus2_4_.oe_async_reset = "none";
defparam ledr_triBus2_4_.oe_power_up = "low";
defparam ledr_triBus2_4_.oe_register_mode = "none";
defparam ledr_triBus2_4_.oe_sync_reset = "none";
defparam ledr_triBus2_4_.operation_mode = "output";
defparam ledr_triBus2_4_.output_async_reset = "none";
defparam ledr_triBus2_4_.output_power_up = "low";
defparam ledr_triBus2_4_.output_register_mode = "none";
defparam ledr_triBus2_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AD23
cycloneii_io ledr_triBus2_5_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[5]));
// synopsys translate_off
defparam ledr_triBus2_5_.input_async_reset = "none";
defparam ledr_triBus2_5_.input_power_up = "low";
defparam ledr_triBus2_5_.input_register_mode = "none";
defparam ledr_triBus2_5_.input_sync_reset = "none";
defparam ledr_triBus2_5_.oe_async_reset = "none";
defparam ledr_triBus2_5_.oe_power_up = "low";
defparam ledr_triBus2_5_.oe_register_mode = "none";
defparam ledr_triBus2_5_.oe_sync_reset = "none";
defparam ledr_triBus2_5_.operation_mode = "output";
defparam ledr_triBus2_5_.output_async_reset = "none";
defparam ledr_triBus2_5_.output_power_up = "low";
defparam ledr_triBus2_5_.output_register_mode = "none";
defparam ledr_triBus2_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AD21
cycloneii_io ledr_triBus2_6_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[6]));
// synopsys translate_off
defparam ledr_triBus2_6_.input_async_reset = "none";
defparam ledr_triBus2_6_.input_power_up = "low";
defparam ledr_triBus2_6_.input_register_mode = "none";
defparam ledr_triBus2_6_.input_sync_reset = "none";
defparam ledr_triBus2_6_.oe_async_reset = "none";
defparam ledr_triBus2_6_.oe_power_up = "low";
defparam ledr_triBus2_6_.oe_register_mode = "none";
defparam ledr_triBus2_6_.oe_sync_reset = "none";
defparam ledr_triBus2_6_.operation_mode = "output";
defparam ledr_triBus2_6_.output_async_reset = "none";
defparam ledr_triBus2_6_.output_power_up = "low";
defparam ledr_triBus2_6_.output_register_mode = "none";
defparam ledr_triBus2_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AC21
cycloneii_io ledr_triBus2_7_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[7]));
// synopsys translate_off
defparam ledr_triBus2_7_.input_async_reset = "none";
defparam ledr_triBus2_7_.input_power_up = "low";
defparam ledr_triBus2_7_.input_register_mode = "none";
defparam ledr_triBus2_7_.input_sync_reset = "none";
defparam ledr_triBus2_7_.oe_async_reset = "none";
defparam ledr_triBus2_7_.oe_power_up = "low";
defparam ledr_triBus2_7_.oe_register_mode = "none";
defparam ledr_triBus2_7_.oe_sync_reset = "none";
defparam ledr_triBus2_7_.operation_mode = "output";
defparam ledr_triBus2_7_.output_async_reset = "none";
defparam ledr_triBus2_7_.output_power_up = "low";
defparam ledr_triBus2_7_.output_register_mode = "none";
defparam ledr_triBus2_7_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AA14
cycloneii_io ledr_triBus2_8_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[8]));
// synopsys translate_off
defparam ledr_triBus2_8_.input_async_reset = "none";
defparam ledr_triBus2_8_.input_power_up = "low";
defparam ledr_triBus2_8_.input_register_mode = "none";
defparam ledr_triBus2_8_.input_sync_reset = "none";
defparam ledr_triBus2_8_.oe_async_reset = "none";
defparam ledr_triBus2_8_.oe_power_up = "low";
defparam ledr_triBus2_8_.oe_register_mode = "none";
defparam ledr_triBus2_8_.oe_sync_reset = "none";
defparam ledr_triBus2_8_.operation_mode = "output";
defparam ledr_triBus2_8_.output_async_reset = "none";
defparam ledr_triBus2_8_.output_power_up = "low";
defparam ledr_triBus2_8_.output_register_mode = "none";
defparam ledr_triBus2_8_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_Y13
cycloneii_io ledr_triBus2_9_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[9]));
// synopsys translate_off
defparam ledr_triBus2_9_.input_async_reset = "none";
defparam ledr_triBus2_9_.input_power_up = "low";
defparam ledr_triBus2_9_.input_register_mode = "none";
defparam ledr_triBus2_9_.input_sync_reset = "none";
defparam ledr_triBus2_9_.oe_async_reset = "none";
defparam ledr_triBus2_9_.oe_power_up = "low";
defparam ledr_triBus2_9_.oe_register_mode = "none";
defparam ledr_triBus2_9_.oe_sync_reset = "none";
defparam ledr_triBus2_9_.operation_mode = "output";
defparam ledr_triBus2_9_.output_async_reset = "none";
defparam ledr_triBus2_9_.output_power_up = "low";
defparam ledr_triBus2_9_.output_register_mode = "none";
defparam ledr_triBus2_9_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AA13
cycloneii_io ledr_triBus2_10_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[10]));
// synopsys translate_off
defparam ledr_triBus2_10_.input_async_reset = "none";
defparam ledr_triBus2_10_.input_power_up = "low";
defparam ledr_triBus2_10_.input_register_mode = "none";
defparam ledr_triBus2_10_.input_sync_reset = "none";
defparam ledr_triBus2_10_.oe_async_reset = "none";
defparam ledr_triBus2_10_.oe_power_up = "low";
defparam ledr_triBus2_10_.oe_register_mode = "none";
defparam ledr_triBus2_10_.oe_sync_reset = "none";
defparam ledr_triBus2_10_.operation_mode = "output";
defparam ledr_triBus2_10_.output_async_reset = "none";
defparam ledr_triBus2_10_.output_power_up = "low";
defparam ledr_triBus2_10_.output_register_mode = "none";
defparam ledr_triBus2_10_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AC14
cycloneii_io ledr_triBus2_11_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[11]));
// synopsys translate_off
defparam ledr_triBus2_11_.input_async_reset = "none";
defparam ledr_triBus2_11_.input_power_up = "low";
defparam ledr_triBus2_11_.input_register_mode = "none";
defparam ledr_triBus2_11_.input_sync_reset = "none";
defparam ledr_triBus2_11_.oe_async_reset = "none";
defparam ledr_triBus2_11_.oe_power_up = "low";
defparam ledr_triBus2_11_.oe_register_mode = "none";
defparam ledr_triBus2_11_.oe_sync_reset = "none";
defparam ledr_triBus2_11_.operation_mode = "output";
defparam ledr_triBus2_11_.output_async_reset = "none";
defparam ledr_triBus2_11_.output_power_up = "low";
defparam ledr_triBus2_11_.output_register_mode = "none";
defparam ledr_triBus2_11_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AD15
cycloneii_io ledr_triBus2_12_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[12]));
// synopsys translate_off
defparam ledr_triBus2_12_.input_async_reset = "none";
defparam ledr_triBus2_12_.input_power_up = "low";
defparam ledr_triBus2_12_.input_register_mode = "none";
defparam ledr_triBus2_12_.input_sync_reset = "none";
defparam ledr_triBus2_12_.oe_async_reset = "none";
defparam ledr_triBus2_12_.oe_power_up = "low";
defparam ledr_triBus2_12_.oe_register_mode = "none";
defparam ledr_triBus2_12_.oe_sync_reset = "none";
defparam ledr_triBus2_12_.operation_mode = "output";
defparam ledr_triBus2_12_.output_async_reset = "none";
defparam ledr_triBus2_12_.output_power_up = "low";
defparam ledr_triBus2_12_.output_register_mode = "none";
defparam ledr_triBus2_12_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AE15
cycloneii_io ledr_triBus2_13_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[13]));
// synopsys translate_off
defparam ledr_triBus2_13_.input_async_reset = "none";
defparam ledr_triBus2_13_.input_power_up = "low";
defparam ledr_triBus2_13_.input_register_mode = "none";
defparam ledr_triBus2_13_.input_sync_reset = "none";
defparam ledr_triBus2_13_.oe_async_reset = "none";
defparam ledr_triBus2_13_.oe_power_up = "low";
defparam ledr_triBus2_13_.oe_register_mode = "none";
defparam ledr_triBus2_13_.oe_sync_reset = "none";
defparam ledr_triBus2_13_.operation_mode = "output";
defparam ledr_triBus2_13_.output_async_reset = "none";
defparam ledr_triBus2_13_.output_power_up = "low";
defparam ledr_triBus2_13_.output_register_mode = "none";
defparam ledr_triBus2_13_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AF13
cycloneii_io ledr_triBus2_14_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[14]));
// synopsys translate_off
defparam ledr_triBus2_14_.input_async_reset = "none";
defparam ledr_triBus2_14_.input_power_up = "low";
defparam ledr_triBus2_14_.input_register_mode = "none";
defparam ledr_triBus2_14_.input_sync_reset = "none";
defparam ledr_triBus2_14_.oe_async_reset = "none";
defparam ledr_triBus2_14_.oe_power_up = "low";
defparam ledr_triBus2_14_.oe_register_mode = "none";
defparam ledr_triBus2_14_.oe_sync_reset = "none";
defparam ledr_triBus2_14_.operation_mode = "output";
defparam ledr_triBus2_14_.output_async_reset = "none";
defparam ledr_triBus2_14_.output_power_up = "low";
defparam ledr_triBus2_14_.output_register_mode = "none";
defparam ledr_triBus2_14_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AE13
cycloneii_io ledr_triBus2_15_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[15]));
// synopsys translate_off
defparam ledr_triBus2_15_.input_async_reset = "none";
defparam ledr_triBus2_15_.input_power_up = "low";
defparam ledr_triBus2_15_.input_register_mode = "none";
defparam ledr_triBus2_15_.input_sync_reset = "none";
defparam ledr_triBus2_15_.oe_async_reset = "none";
defparam ledr_triBus2_15_.oe_power_up = "low";
defparam ledr_triBus2_15_.oe_register_mode = "none";
defparam ledr_triBus2_15_.oe_sync_reset = "none";
defparam ledr_triBus2_15_.operation_mode = "output";
defparam ledr_triBus2_15_.output_async_reset = "none";
defparam ledr_triBus2_15_.output_power_up = "low";
defparam ledr_triBus2_15_.output_register_mode = "none";
defparam ledr_triBus2_15_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AE12
cycloneii_io ledr_triBus2_16_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[16]));
// synopsys translate_off
defparam ledr_triBus2_16_.input_async_reset = "none";
defparam ledr_triBus2_16_.input_power_up = "low";
defparam ledr_triBus2_16_.input_register_mode = "none";
defparam ledr_triBus2_16_.input_sync_reset = "none";
defparam ledr_triBus2_16_.oe_async_reset = "none";
defparam ledr_triBus2_16_.oe_power_up = "low";
defparam ledr_triBus2_16_.oe_register_mode = "none";
defparam ledr_triBus2_16_.oe_sync_reset = "none";
defparam ledr_triBus2_16_.operation_mode = "output";
defparam ledr_triBus2_16_.output_async_reset = "none";
defparam ledr_triBus2_16_.output_power_up = "low";
defparam ledr_triBus2_16_.output_register_mode = "none";
defparam ledr_triBus2_16_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AD12
cycloneii_io ledr_triBus2_17_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(ledr[17]));
// synopsys translate_off
defparam ledr_triBus2_17_.input_async_reset = "none";
defparam ledr_triBus2_17_.input_power_up = "low";
defparam ledr_triBus2_17_.input_register_mode = "none";
defparam ledr_triBus2_17_.input_sync_reset = "none";
defparam ledr_triBus2_17_.oe_async_reset = "none";
defparam ledr_triBus2_17_.oe_power_up = "low";
defparam ledr_triBus2_17_.oe_register_mode = "none";
defparam ledr_triBus2_17_.oe_sync_reset = "none";
defparam ledr_triBus2_17_.operation_mode = "output";
defparam ledr_triBus2_17_.output_async_reset = "none";
defparam ledr_triBus2_17_.output_power_up = "low";
defparam ledr_triBus2_17_.output_register_mode = "none";
defparam ledr_triBus2_17_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AF10
cycloneii_io hex0_triBus3_0_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex0[0]));
// synopsys translate_off
defparam hex0_triBus3_0_.input_async_reset = "none";
defparam hex0_triBus3_0_.input_power_up = "low";
defparam hex0_triBus3_0_.input_register_mode = "none";
defparam hex0_triBus3_0_.input_sync_reset = "none";
defparam hex0_triBus3_0_.oe_async_reset = "none";
defparam hex0_triBus3_0_.oe_power_up = "low";
defparam hex0_triBus3_0_.oe_register_mode = "none";
defparam hex0_triBus3_0_.oe_sync_reset = "none";
defparam hex0_triBus3_0_.operation_mode = "output";
defparam hex0_triBus3_0_.output_async_reset = "none";
defparam hex0_triBus3_0_.output_power_up = "low";
defparam hex0_triBus3_0_.output_register_mode = "none";
defparam hex0_triBus3_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AB12
cycloneii_io hex0_triBus3_1_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex0[1]));
// synopsys translate_off
defparam hex0_triBus3_1_.input_async_reset = "none";
defparam hex0_triBus3_1_.input_power_up = "low";
defparam hex0_triBus3_1_.input_register_mode = "none";
defparam hex0_triBus3_1_.input_sync_reset = "none";
defparam hex0_triBus3_1_.oe_async_reset = "none";
defparam hex0_triBus3_1_.oe_power_up = "low";
defparam hex0_triBus3_1_.oe_register_mode = "none";
defparam hex0_triBus3_1_.oe_sync_reset = "none";
defparam hex0_triBus3_1_.operation_mode = "output";
defparam hex0_triBus3_1_.output_async_reset = "none";
defparam hex0_triBus3_1_.output_power_up = "low";
defparam hex0_triBus3_1_.output_register_mode = "none";
defparam hex0_triBus3_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AC12
cycloneii_io hex0_triBus3_2_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex0[2]));
// synopsys translate_off
defparam hex0_triBus3_2_.input_async_reset = "none";
defparam hex0_triBus3_2_.input_power_up = "low";
defparam hex0_triBus3_2_.input_register_mode = "none";
defparam hex0_triBus3_2_.input_sync_reset = "none";
defparam hex0_triBus3_2_.oe_async_reset = "none";
defparam hex0_triBus3_2_.oe_power_up = "low";
defparam hex0_triBus3_2_.oe_register_mode = "none";
defparam hex0_triBus3_2_.oe_sync_reset = "none";
defparam hex0_triBus3_2_.operation_mode = "output";
defparam hex0_triBus3_2_.output_async_reset = "none";
defparam hex0_triBus3_2_.output_power_up = "low";
defparam hex0_triBus3_2_.output_register_mode = "none";
defparam hex0_triBus3_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AD11
cycloneii_io hex0_triBus3_3_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex0[3]));
// synopsys translate_off
defparam hex0_triBus3_3_.input_async_reset = "none";
defparam hex0_triBus3_3_.input_power_up = "low";
defparam hex0_triBus3_3_.input_register_mode = "none";
defparam hex0_triBus3_3_.input_sync_reset = "none";
defparam hex0_triBus3_3_.oe_async_reset = "none";
defparam hex0_triBus3_3_.oe_power_up = "low";
defparam hex0_triBus3_3_.oe_register_mode = "none";
defparam hex0_triBus3_3_.oe_sync_reset = "none";
defparam hex0_triBus3_3_.operation_mode = "output";
defparam hex0_triBus3_3_.output_async_reset = "none";
defparam hex0_triBus3_3_.output_power_up = "low";
defparam hex0_triBus3_3_.output_register_mode = "none";
defparam hex0_triBus3_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AE11
cycloneii_io hex0_triBus3_4_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex0[4]));
// synopsys translate_off
defparam hex0_triBus3_4_.input_async_reset = "none";
defparam hex0_triBus3_4_.input_power_up = "low";
defparam hex0_triBus3_4_.input_register_mode = "none";
defparam hex0_triBus3_4_.input_sync_reset = "none";
defparam hex0_triBus3_4_.oe_async_reset = "none";
defparam hex0_triBus3_4_.oe_power_up = "low";
defparam hex0_triBus3_4_.oe_register_mode = "none";
defparam hex0_triBus3_4_.oe_sync_reset = "none";
defparam hex0_triBus3_4_.operation_mode = "output";
defparam hex0_triBus3_4_.output_async_reset = "none";
defparam hex0_triBus3_4_.output_power_up = "low";
defparam hex0_triBus3_4_.output_register_mode = "none";
defparam hex0_triBus3_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_V14
cycloneii_io hex0_triBus3_5_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex0[5]));
// synopsys translate_off
defparam hex0_triBus3_5_.input_async_reset = "none";
defparam hex0_triBus3_5_.input_power_up = "low";
defparam hex0_triBus3_5_.input_register_mode = "none";
defparam hex0_triBus3_5_.input_sync_reset = "none";
defparam hex0_triBus3_5_.oe_async_reset = "none";
defparam hex0_triBus3_5_.oe_power_up = "low";
defparam hex0_triBus3_5_.oe_register_mode = "none";
defparam hex0_triBus3_5_.oe_sync_reset = "none";
defparam hex0_triBus3_5_.operation_mode = "output";
defparam hex0_triBus3_5_.output_async_reset = "none";
defparam hex0_triBus3_5_.output_power_up = "low";
defparam hex0_triBus3_5_.output_register_mode = "none";
defparam hex0_triBus3_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_V13
cycloneii_io hex0_triBus3_6_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex0[6]));
// synopsys translate_off
defparam hex0_triBus3_6_.input_async_reset = "none";
defparam hex0_triBus3_6_.input_power_up = "low";
defparam hex0_triBus3_6_.input_register_mode = "none";
defparam hex0_triBus3_6_.input_sync_reset = "none";
defparam hex0_triBus3_6_.oe_async_reset = "none";
defparam hex0_triBus3_6_.oe_power_up = "low";
defparam hex0_triBus3_6_.oe_register_mode = "none";
defparam hex0_triBus3_6_.oe_sync_reset = "none";
defparam hex0_triBus3_6_.operation_mode = "output";
defparam hex0_triBus3_6_.output_async_reset = "none";
defparam hex0_triBus3_6_.output_power_up = "low";
defparam hex0_triBus3_6_.output_register_mode = "none";
defparam hex0_triBus3_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_V20
cycloneii_io hex1_triBus4_0_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex1[0]));
// synopsys translate_off
defparam hex1_triBus4_0_.input_async_reset = "none";
defparam hex1_triBus4_0_.input_power_up = "low";
defparam hex1_triBus4_0_.input_register_mode = "none";
defparam hex1_triBus4_0_.input_sync_reset = "none";
defparam hex1_triBus4_0_.oe_async_reset = "none";
defparam hex1_triBus4_0_.oe_power_up = "low";
defparam hex1_triBus4_0_.oe_register_mode = "none";
defparam hex1_triBus4_0_.oe_sync_reset = "none";
defparam hex1_triBus4_0_.operation_mode = "output";
defparam hex1_triBus4_0_.output_async_reset = "none";
defparam hex1_triBus4_0_.output_power_up = "low";
defparam hex1_triBus4_0_.output_register_mode = "none";
defparam hex1_triBus4_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_V21
cycloneii_io hex1_triBus4_1_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex1[1]));
// synopsys translate_off
defparam hex1_triBus4_1_.input_async_reset = "none";
defparam hex1_triBus4_1_.input_power_up = "low";
defparam hex1_triBus4_1_.input_register_mode = "none";
defparam hex1_triBus4_1_.input_sync_reset = "none";
defparam hex1_triBus4_1_.oe_async_reset = "none";
defparam hex1_triBus4_1_.oe_power_up = "low";
defparam hex1_triBus4_1_.oe_register_mode = "none";
defparam hex1_triBus4_1_.oe_sync_reset = "none";
defparam hex1_triBus4_1_.operation_mode = "output";
defparam hex1_triBus4_1_.output_async_reset = "none";
defparam hex1_triBus4_1_.output_power_up = "low";
defparam hex1_triBus4_1_.output_register_mode = "none";
defparam hex1_triBus4_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_W21
cycloneii_io hex1_triBus4_2_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex1[2]));
// synopsys translate_off
defparam hex1_triBus4_2_.input_async_reset = "none";
defparam hex1_triBus4_2_.input_power_up = "low";
defparam hex1_triBus4_2_.input_register_mode = "none";
defparam hex1_triBus4_2_.input_sync_reset = "none";
defparam hex1_triBus4_2_.oe_async_reset = "none";
defparam hex1_triBus4_2_.oe_power_up = "low";
defparam hex1_triBus4_2_.oe_register_mode = "none";
defparam hex1_triBus4_2_.oe_sync_reset = "none";
defparam hex1_triBus4_2_.operation_mode = "output";
defparam hex1_triBus4_2_.output_async_reset = "none";
defparam hex1_triBus4_2_.output_power_up = "low";
defparam hex1_triBus4_2_.output_register_mode = "none";
defparam hex1_triBus4_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_Y22
cycloneii_io hex1_triBus4_3_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex1[3]));
// synopsys translate_off
defparam hex1_triBus4_3_.input_async_reset = "none";
defparam hex1_triBus4_3_.input_power_up = "low";
defparam hex1_triBus4_3_.input_register_mode = "none";
defparam hex1_triBus4_3_.input_sync_reset = "none";
defparam hex1_triBus4_3_.oe_async_reset = "none";
defparam hex1_triBus4_3_.oe_power_up = "low";
defparam hex1_triBus4_3_.oe_register_mode = "none";
defparam hex1_triBus4_3_.oe_sync_reset = "none";
defparam hex1_triBus4_3_.operation_mode = "output";
defparam hex1_triBus4_3_.output_async_reset = "none";
defparam hex1_triBus4_3_.output_power_up = "low";
defparam hex1_triBus4_3_.output_register_mode = "none";
defparam hex1_triBus4_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AA24
cycloneii_io hex1_triBus4_4_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex1[4]));
// synopsys translate_off
defparam hex1_triBus4_4_.input_async_reset = "none";
defparam hex1_triBus4_4_.input_power_up = "low";
defparam hex1_triBus4_4_.input_register_mode = "none";
defparam hex1_triBus4_4_.input_sync_reset = "none";
defparam hex1_triBus4_4_.oe_async_reset = "none";
defparam hex1_triBus4_4_.oe_power_up = "low";
defparam hex1_triBus4_4_.oe_register_mode = "none";
defparam hex1_triBus4_4_.oe_sync_reset = "none";
defparam hex1_triBus4_4_.operation_mode = "output";
defparam hex1_triBus4_4_.output_async_reset = "none";
defparam hex1_triBus4_4_.output_power_up = "low";
defparam hex1_triBus4_4_.output_register_mode = "none";
defparam hex1_triBus4_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AA23
cycloneii_io hex1_triBus4_5_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex1[5]));
// synopsys translate_off
defparam hex1_triBus4_5_.input_async_reset = "none";
defparam hex1_triBus4_5_.input_power_up = "low";
defparam hex1_triBus4_5_.input_register_mode = "none";
defparam hex1_triBus4_5_.input_sync_reset = "none";
defparam hex1_triBus4_5_.oe_async_reset = "none";
defparam hex1_triBus4_5_.oe_power_up = "low";
defparam hex1_triBus4_5_.oe_register_mode = "none";
defparam hex1_triBus4_5_.oe_sync_reset = "none";
defparam hex1_triBus4_5_.operation_mode = "output";
defparam hex1_triBus4_5_.output_async_reset = "none";
defparam hex1_triBus4_5_.output_power_up = "low";
defparam hex1_triBus4_5_.output_register_mode = "none";
defparam hex1_triBus4_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AB24
cycloneii_io hex1_triBus4_6_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex1[6]));
// synopsys translate_off
defparam hex1_triBus4_6_.input_async_reset = "none";
defparam hex1_triBus4_6_.input_power_up = "low";
defparam hex1_triBus4_6_.input_register_mode = "none";
defparam hex1_triBus4_6_.input_sync_reset = "none";
defparam hex1_triBus4_6_.oe_async_reset = "none";
defparam hex1_triBus4_6_.oe_power_up = "low";
defparam hex1_triBus4_6_.oe_register_mode = "none";
defparam hex1_triBus4_6_.oe_sync_reset = "none";
defparam hex1_triBus4_6_.operation_mode = "output";
defparam hex1_triBus4_6_.output_async_reset = "none";
defparam hex1_triBus4_6_.output_power_up = "low";
defparam hex1_triBus4_6_.output_register_mode = "none";
defparam hex1_triBus4_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AB23
cycloneii_io hex2_triBus5_0_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex2[0]));
// synopsys translate_off
defparam hex2_triBus5_0_.input_async_reset = "none";
defparam hex2_triBus5_0_.input_power_up = "low";
defparam hex2_triBus5_0_.input_register_mode = "none";
defparam hex2_triBus5_0_.input_sync_reset = "none";
defparam hex2_triBus5_0_.oe_async_reset = "none";
defparam hex2_triBus5_0_.oe_power_up = "low";
defparam hex2_triBus5_0_.oe_register_mode = "none";
defparam hex2_triBus5_0_.oe_sync_reset = "none";
defparam hex2_triBus5_0_.operation_mode = "output";
defparam hex2_triBus5_0_.output_async_reset = "none";
defparam hex2_triBus5_0_.output_power_up = "low";
defparam hex2_triBus5_0_.output_register_mode = "none";
defparam hex2_triBus5_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_V22
cycloneii_io hex2_triBus5_1_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex2[1]));
// synopsys translate_off
defparam hex2_triBus5_1_.input_async_reset = "none";
defparam hex2_triBus5_1_.input_power_up = "low";
defparam hex2_triBus5_1_.input_register_mode = "none";
defparam hex2_triBus5_1_.input_sync_reset = "none";
defparam hex2_triBus5_1_.oe_async_reset = "none";
defparam hex2_triBus5_1_.oe_power_up = "low";
defparam hex2_triBus5_1_.oe_register_mode = "none";
defparam hex2_triBus5_1_.oe_sync_reset = "none";
defparam hex2_triBus5_1_.operation_mode = "output";
defparam hex2_triBus5_1_.output_async_reset = "none";
defparam hex2_triBus5_1_.output_power_up = "low";
defparam hex2_triBus5_1_.output_register_mode = "none";
defparam hex2_triBus5_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AC25
cycloneii_io hex2_triBus5_2_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex2[2]));
// synopsys translate_off
defparam hex2_triBus5_2_.input_async_reset = "none";
defparam hex2_triBus5_2_.input_power_up = "low";
defparam hex2_triBus5_2_.input_register_mode = "none";
defparam hex2_triBus5_2_.input_sync_reset = "none";
defparam hex2_triBus5_2_.oe_async_reset = "none";
defparam hex2_triBus5_2_.oe_power_up = "low";
defparam hex2_triBus5_2_.oe_register_mode = "none";
defparam hex2_triBus5_2_.oe_sync_reset = "none";
defparam hex2_triBus5_2_.operation_mode = "output";
defparam hex2_triBus5_2_.output_async_reset = "none";
defparam hex2_triBus5_2_.output_power_up = "low";
defparam hex2_triBus5_2_.output_register_mode = "none";
defparam hex2_triBus5_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AC26
cycloneii_io hex2_triBus5_3_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex2[3]));
// synopsys translate_off
defparam hex2_triBus5_3_.input_async_reset = "none";
defparam hex2_triBus5_3_.input_power_up = "low";
defparam hex2_triBus5_3_.input_register_mode = "none";
defparam hex2_triBus5_3_.input_sync_reset = "none";
defparam hex2_triBus5_3_.oe_async_reset = "none";
defparam hex2_triBus5_3_.oe_power_up = "low";
defparam hex2_triBus5_3_.oe_register_mode = "none";
defparam hex2_triBus5_3_.oe_sync_reset = "none";
defparam hex2_triBus5_3_.operation_mode = "output";
defparam hex2_triBus5_3_.output_async_reset = "none";
defparam hex2_triBus5_3_.output_power_up = "low";
defparam hex2_triBus5_3_.output_register_mode = "none";
defparam hex2_triBus5_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AB26
cycloneii_io hex2_triBus5_4_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex2[4]));
// synopsys translate_off
defparam hex2_triBus5_4_.input_async_reset = "none";
defparam hex2_triBus5_4_.input_power_up = "low";
defparam hex2_triBus5_4_.input_register_mode = "none";
defparam hex2_triBus5_4_.input_sync_reset = "none";
defparam hex2_triBus5_4_.oe_async_reset = "none";
defparam hex2_triBus5_4_.oe_power_up = "low";
defparam hex2_triBus5_4_.oe_register_mode = "none";
defparam hex2_triBus5_4_.oe_sync_reset = "none";
defparam hex2_triBus5_4_.operation_mode = "output";
defparam hex2_triBus5_4_.output_async_reset = "none";
defparam hex2_triBus5_4_.output_power_up = "low";
defparam hex2_triBus5_4_.output_register_mode = "none";
defparam hex2_triBus5_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AB25
cycloneii_io hex2_triBus5_5_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex2[5]));
// synopsys translate_off
defparam hex2_triBus5_5_.input_async_reset = "none";
defparam hex2_triBus5_5_.input_power_up = "low";
defparam hex2_triBus5_5_.input_register_mode = "none";
defparam hex2_triBus5_5_.input_sync_reset = "none";
defparam hex2_triBus5_5_.oe_async_reset = "none";
defparam hex2_triBus5_5_.oe_power_up = "low";
defparam hex2_triBus5_5_.oe_register_mode = "none";
defparam hex2_triBus5_5_.oe_sync_reset = "none";
defparam hex2_triBus5_5_.operation_mode = "output";
defparam hex2_triBus5_5_.output_async_reset = "none";
defparam hex2_triBus5_5_.output_power_up = "low";
defparam hex2_triBus5_5_.output_register_mode = "none";
defparam hex2_triBus5_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_Y24
cycloneii_io hex2_triBus5_6_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex2[6]));
// synopsys translate_off
defparam hex2_triBus5_6_.input_async_reset = "none";
defparam hex2_triBus5_6_.input_power_up = "low";
defparam hex2_triBus5_6_.input_register_mode = "none";
defparam hex2_triBus5_6_.input_sync_reset = "none";
defparam hex2_triBus5_6_.oe_async_reset = "none";
defparam hex2_triBus5_6_.oe_power_up = "low";
defparam hex2_triBus5_6_.oe_register_mode = "none";
defparam hex2_triBus5_6_.oe_sync_reset = "none";
defparam hex2_triBus5_6_.operation_mode = "output";
defparam hex2_triBus5_6_.output_async_reset = "none";
defparam hex2_triBus5_6_.output_power_up = "low";
defparam hex2_triBus5_6_.output_register_mode = "none";
defparam hex2_triBus5_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_Y23
cycloneii_io hex3_triBus6_0_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex3[0]));
// synopsys translate_off
defparam hex3_triBus6_0_.input_async_reset = "none";
defparam hex3_triBus6_0_.input_power_up = "low";
defparam hex3_triBus6_0_.input_register_mode = "none";
defparam hex3_triBus6_0_.input_sync_reset = "none";
defparam hex3_triBus6_0_.oe_async_reset = "none";
defparam hex3_triBus6_0_.oe_power_up = "low";
defparam hex3_triBus6_0_.oe_register_mode = "none";
defparam hex3_triBus6_0_.oe_sync_reset = "none";
defparam hex3_triBus6_0_.operation_mode = "output";
defparam hex3_triBus6_0_.output_async_reset = "none";
defparam hex3_triBus6_0_.output_power_up = "low";
defparam hex3_triBus6_0_.output_register_mode = "none";
defparam hex3_triBus6_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AA25
cycloneii_io hex3_triBus6_1_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex3[1]));
// synopsys translate_off
defparam hex3_triBus6_1_.input_async_reset = "none";
defparam hex3_triBus6_1_.input_power_up = "low";
defparam hex3_triBus6_1_.input_register_mode = "none";
defparam hex3_triBus6_1_.input_sync_reset = "none";
defparam hex3_triBus6_1_.oe_async_reset = "none";
defparam hex3_triBus6_1_.oe_power_up = "low";
defparam hex3_triBus6_1_.oe_register_mode = "none";
defparam hex3_triBus6_1_.oe_sync_reset = "none";
defparam hex3_triBus6_1_.operation_mode = "output";
defparam hex3_triBus6_1_.output_async_reset = "none";
defparam hex3_triBus6_1_.output_power_up = "low";
defparam hex3_triBus6_1_.output_register_mode = "none";
defparam hex3_triBus6_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_AA26
cycloneii_io hex3_triBus6_2_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex3[2]));
// synopsys translate_off
defparam hex3_triBus6_2_.input_async_reset = "none";
defparam hex3_triBus6_2_.input_power_up = "low";
defparam hex3_triBus6_2_.input_register_mode = "none";
defparam hex3_triBus6_2_.input_sync_reset = "none";
defparam hex3_triBus6_2_.oe_async_reset = "none";
defparam hex3_triBus6_2_.oe_power_up = "low";
defparam hex3_triBus6_2_.oe_register_mode = "none";
defparam hex3_triBus6_2_.oe_sync_reset = "none";
defparam hex3_triBus6_2_.operation_mode = "output";
defparam hex3_triBus6_2_.output_async_reset = "none";
defparam hex3_triBus6_2_.output_power_up = "low";
defparam hex3_triBus6_2_.output_register_mode = "none";
defparam hex3_triBus6_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_Y26
cycloneii_io hex3_triBus6_3_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex3[3]));
// synopsys translate_off
defparam hex3_triBus6_3_.input_async_reset = "none";
defparam hex3_triBus6_3_.input_power_up = "low";
defparam hex3_triBus6_3_.input_register_mode = "none";
defparam hex3_triBus6_3_.input_sync_reset = "none";
defparam hex3_triBus6_3_.oe_async_reset = "none";
defparam hex3_triBus6_3_.oe_power_up = "low";
defparam hex3_triBus6_3_.oe_register_mode = "none";
defparam hex3_triBus6_3_.oe_sync_reset = "none";
defparam hex3_triBus6_3_.operation_mode = "output";
defparam hex3_triBus6_3_.output_async_reset = "none";
defparam hex3_triBus6_3_.output_power_up = "low";
defparam hex3_triBus6_3_.output_register_mode = "none";
defparam hex3_triBus6_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_Y25
cycloneii_io hex3_triBus6_4_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex3[4]));
// synopsys translate_off
defparam hex3_triBus6_4_.input_async_reset = "none";
defparam hex3_triBus6_4_.input_power_up = "low";
defparam hex3_triBus6_4_.input_register_mode = "none";
defparam hex3_triBus6_4_.input_sync_reset = "none";
defparam hex3_triBus6_4_.oe_async_reset = "none";
defparam hex3_triBus6_4_.oe_power_up = "low";
defparam hex3_triBus6_4_.oe_register_mode = "none";
defparam hex3_triBus6_4_.oe_sync_reset = "none";
defparam hex3_triBus6_4_.operation_mode = "output";
defparam hex3_triBus6_4_.output_async_reset = "none";
defparam hex3_triBus6_4_.output_power_up = "low";
defparam hex3_triBus6_4_.output_register_mode = "none";
defparam hex3_triBus6_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_U22
cycloneii_io hex3_triBus6_5_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex3[5]));
// synopsys translate_off
defparam hex3_triBus6_5_.input_async_reset = "none";
defparam hex3_triBus6_5_.input_power_up = "low";
defparam hex3_triBus6_5_.input_register_mode = "none";
defparam hex3_triBus6_5_.input_sync_reset = "none";
defparam hex3_triBus6_5_.oe_async_reset = "none";
defparam hex3_triBus6_5_.oe_power_up = "low";
defparam hex3_triBus6_5_.oe_register_mode = "none";
defparam hex3_triBus6_5_.oe_sync_reset = "none";
defparam hex3_triBus6_5_.operation_mode = "output";
defparam hex3_triBus6_5_.output_async_reset = "none";
defparam hex3_triBus6_5_.output_power_up = "low";
defparam hex3_triBus6_5_.output_register_mode = "none";
defparam hex3_triBus6_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_W24
cycloneii_io hex3_triBus6_6_(
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex3[6]));
// synopsys translate_off
defparam hex3_triBus6_6_.input_async_reset = "none";
defparam hex3_triBus6_6_.input_power_up = "low";
defparam hex3_triBus6_6_.input_register_mode = "none";
defparam hex3_triBus6_6_.input_sync_reset = "none";
defparam hex3_triBus6_6_.oe_async_reset = "none";
defparam hex3_triBus6_6_.oe_power_up = "low";
defparam hex3_triBus6_6_.oe_register_mode = "none";
defparam hex3_triBus6_6_.oe_sync_reset = "none";
defparam hex3_triBus6_6_.operation_mode = "output";
defparam hex3_triBus6_6_.output_async_reset = "none";
defparam hex3_triBus6_6_.output_power_up = "low";
defparam hex3_triBus6_6_.output_register_mode = "none";
defparam hex3_triBus6_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_U9
cycloneii_io hex4_obuf_0_(
	.datain(hex4_dup0_0_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex4[0]));
// synopsys translate_off
defparam hex4_obuf_0_.input_async_reset = "none";
defparam hex4_obuf_0_.input_power_up = "low";
defparam hex4_obuf_0_.input_register_mode = "none";
defparam hex4_obuf_0_.input_sync_reset = "none";
defparam hex4_obuf_0_.oe_async_reset = "none";
defparam hex4_obuf_0_.oe_power_up = "low";
defparam hex4_obuf_0_.oe_register_mode = "none";
defparam hex4_obuf_0_.oe_sync_reset = "none";
defparam hex4_obuf_0_.operation_mode = "output";
defparam hex4_obuf_0_.output_async_reset = "none";
defparam hex4_obuf_0_.output_power_up = "low";
defparam hex4_obuf_0_.output_register_mode = "none";
defparam hex4_obuf_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_U1
cycloneii_io hex4_obuf_1_(
	.datain(hex4_dup0_1_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex4[1]));
// synopsys translate_off
defparam hex4_obuf_1_.input_async_reset = "none";
defparam hex4_obuf_1_.input_power_up = "low";
defparam hex4_obuf_1_.input_register_mode = "none";
defparam hex4_obuf_1_.input_sync_reset = "none";
defparam hex4_obuf_1_.oe_async_reset = "none";
defparam hex4_obuf_1_.oe_power_up = "low";
defparam hex4_obuf_1_.oe_register_mode = "none";
defparam hex4_obuf_1_.oe_sync_reset = "none";
defparam hex4_obuf_1_.operation_mode = "output";
defparam hex4_obuf_1_.output_async_reset = "none";
defparam hex4_obuf_1_.output_power_up = "low";
defparam hex4_obuf_1_.output_register_mode = "none";
defparam hex4_obuf_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_U2
cycloneii_io hex4_obuf_2_(
	.datain(hex4_dup0_2_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex4[2]));
// synopsys translate_off
defparam hex4_obuf_2_.input_async_reset = "none";
defparam hex4_obuf_2_.input_power_up = "low";
defparam hex4_obuf_2_.input_register_mode = "none";
defparam hex4_obuf_2_.input_sync_reset = "none";
defparam hex4_obuf_2_.oe_async_reset = "none";
defparam hex4_obuf_2_.oe_power_up = "low";
defparam hex4_obuf_2_.oe_register_mode = "none";
defparam hex4_obuf_2_.oe_sync_reset = "none";
defparam hex4_obuf_2_.operation_mode = "output";
defparam hex4_obuf_2_.output_async_reset = "none";
defparam hex4_obuf_2_.output_power_up = "low";
defparam hex4_obuf_2_.output_register_mode = "none";
defparam hex4_obuf_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_T4
cycloneii_io hex4_obuf_3_(
	.datain(hex4_dup0_3_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex4[3]));
// synopsys translate_off
defparam hex4_obuf_3_.input_async_reset = "none";
defparam hex4_obuf_3_.input_power_up = "low";
defparam hex4_obuf_3_.input_register_mode = "none";
defparam hex4_obuf_3_.input_sync_reset = "none";
defparam hex4_obuf_3_.oe_async_reset = "none";
defparam hex4_obuf_3_.oe_power_up = "low";
defparam hex4_obuf_3_.oe_register_mode = "none";
defparam hex4_obuf_3_.oe_sync_reset = "none";
defparam hex4_obuf_3_.operation_mode = "output";
defparam hex4_obuf_3_.output_async_reset = "none";
defparam hex4_obuf_3_.output_power_up = "low";
defparam hex4_obuf_3_.output_register_mode = "none";
defparam hex4_obuf_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_R7
cycloneii_io hex4_obuf_4_(
	.datain(hex4_dup0_4_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex4[4]));
// synopsys translate_off
defparam hex4_obuf_4_.input_async_reset = "none";
defparam hex4_obuf_4_.input_power_up = "low";
defparam hex4_obuf_4_.input_register_mode = "none";
defparam hex4_obuf_4_.input_sync_reset = "none";
defparam hex4_obuf_4_.oe_async_reset = "none";
defparam hex4_obuf_4_.oe_power_up = "low";
defparam hex4_obuf_4_.oe_register_mode = "none";
defparam hex4_obuf_4_.oe_sync_reset = "none";
defparam hex4_obuf_4_.operation_mode = "output";
defparam hex4_obuf_4_.output_async_reset = "none";
defparam hex4_obuf_4_.output_power_up = "low";
defparam hex4_obuf_4_.output_register_mode = "none";
defparam hex4_obuf_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_R6
cycloneii_io hex4_obuf_5_(
	.datain(hex4_dup0_5_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex4[5]));
// synopsys translate_off
defparam hex4_obuf_5_.input_async_reset = "none";
defparam hex4_obuf_5_.input_power_up = "low";
defparam hex4_obuf_5_.input_register_mode = "none";
defparam hex4_obuf_5_.input_sync_reset = "none";
defparam hex4_obuf_5_.oe_async_reset = "none";
defparam hex4_obuf_5_.oe_power_up = "low";
defparam hex4_obuf_5_.oe_register_mode = "none";
defparam hex4_obuf_5_.oe_sync_reset = "none";
defparam hex4_obuf_5_.operation_mode = "output";
defparam hex4_obuf_5_.output_async_reset = "none";
defparam hex4_obuf_5_.output_power_up = "low";
defparam hex4_obuf_5_.output_register_mode = "none";
defparam hex4_obuf_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_T3
cycloneii_io hex4_obuf_6_(
	.datain(hex4_dup0_6_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex4[6]));
// synopsys translate_off
defparam hex4_obuf_6_.input_async_reset = "none";
defparam hex4_obuf_6_.input_power_up = "low";
defparam hex4_obuf_6_.input_register_mode = "none";
defparam hex4_obuf_6_.input_sync_reset = "none";
defparam hex4_obuf_6_.oe_async_reset = "none";
defparam hex4_obuf_6_.oe_power_up = "low";
defparam hex4_obuf_6_.oe_register_mode = "none";
defparam hex4_obuf_6_.oe_sync_reset = "none";
defparam hex4_obuf_6_.operation_mode = "output";
defparam hex4_obuf_6_.output_async_reset = "none";
defparam hex4_obuf_6_.output_power_up = "low";
defparam hex4_obuf_6_.output_register_mode = "none";
defparam hex4_obuf_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_T2
cycloneii_io hex5_obuf_0_(
	.datain(hex5_dup0_0_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex5[0]));
// synopsys translate_off
defparam hex5_obuf_0_.input_async_reset = "none";
defparam hex5_obuf_0_.input_power_up = "low";
defparam hex5_obuf_0_.input_register_mode = "none";
defparam hex5_obuf_0_.input_sync_reset = "none";
defparam hex5_obuf_0_.oe_async_reset = "none";
defparam hex5_obuf_0_.oe_power_up = "low";
defparam hex5_obuf_0_.oe_register_mode = "none";
defparam hex5_obuf_0_.oe_sync_reset = "none";
defparam hex5_obuf_0_.operation_mode = "output";
defparam hex5_obuf_0_.output_async_reset = "none";
defparam hex5_obuf_0_.output_power_up = "low";
defparam hex5_obuf_0_.output_register_mode = "none";
defparam hex5_obuf_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P6
cycloneii_io hex5_obuf_1_(
	.datain(hex5_dup0_1_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex5[1]));
// synopsys translate_off
defparam hex5_obuf_1_.input_async_reset = "none";
defparam hex5_obuf_1_.input_power_up = "low";
defparam hex5_obuf_1_.input_register_mode = "none";
defparam hex5_obuf_1_.input_sync_reset = "none";
defparam hex5_obuf_1_.oe_async_reset = "none";
defparam hex5_obuf_1_.oe_power_up = "low";
defparam hex5_obuf_1_.oe_register_mode = "none";
defparam hex5_obuf_1_.oe_sync_reset = "none";
defparam hex5_obuf_1_.operation_mode = "output";
defparam hex5_obuf_1_.output_async_reset = "none";
defparam hex5_obuf_1_.output_power_up = "low";
defparam hex5_obuf_1_.output_register_mode = "none";
defparam hex5_obuf_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P7
cycloneii_io hex5_obuf_2_(
	.datain(hex5_dup0_2_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex5[2]));
// synopsys translate_off
defparam hex5_obuf_2_.input_async_reset = "none";
defparam hex5_obuf_2_.input_power_up = "low";
defparam hex5_obuf_2_.input_register_mode = "none";
defparam hex5_obuf_2_.input_sync_reset = "none";
defparam hex5_obuf_2_.oe_async_reset = "none";
defparam hex5_obuf_2_.oe_power_up = "low";
defparam hex5_obuf_2_.oe_register_mode = "none";
defparam hex5_obuf_2_.oe_sync_reset = "none";
defparam hex5_obuf_2_.operation_mode = "output";
defparam hex5_obuf_2_.output_async_reset = "none";
defparam hex5_obuf_2_.output_power_up = "low";
defparam hex5_obuf_2_.output_register_mode = "none";
defparam hex5_obuf_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_T9
cycloneii_io hex5_obuf_3_(
	.datain(hex5_dup0_3_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex5[3]));
// synopsys translate_off
defparam hex5_obuf_3_.input_async_reset = "none";
defparam hex5_obuf_3_.input_power_up = "low";
defparam hex5_obuf_3_.input_register_mode = "none";
defparam hex5_obuf_3_.input_sync_reset = "none";
defparam hex5_obuf_3_.oe_async_reset = "none";
defparam hex5_obuf_3_.oe_power_up = "low";
defparam hex5_obuf_3_.oe_register_mode = "none";
defparam hex5_obuf_3_.oe_sync_reset = "none";
defparam hex5_obuf_3_.operation_mode = "output";
defparam hex5_obuf_3_.output_async_reset = "none";
defparam hex5_obuf_3_.output_power_up = "low";
defparam hex5_obuf_3_.output_register_mode = "none";
defparam hex5_obuf_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_R5
cycloneii_io hex5_obuf_4_(
	.datain(hex5_dup0_4_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex5[4]));
// synopsys translate_off
defparam hex5_obuf_4_.input_async_reset = "none";
defparam hex5_obuf_4_.input_power_up = "low";
defparam hex5_obuf_4_.input_register_mode = "none";
defparam hex5_obuf_4_.input_sync_reset = "none";
defparam hex5_obuf_4_.oe_async_reset = "none";
defparam hex5_obuf_4_.oe_power_up = "low";
defparam hex5_obuf_4_.oe_register_mode = "none";
defparam hex5_obuf_4_.oe_sync_reset = "none";
defparam hex5_obuf_4_.operation_mode = "output";
defparam hex5_obuf_4_.output_async_reset = "none";
defparam hex5_obuf_4_.output_power_up = "low";
defparam hex5_obuf_4_.output_register_mode = "none";
defparam hex5_obuf_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_R4
cycloneii_io hex5_obuf_5_(
	.datain(hex5_dup0_5_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex5[5]));
// synopsys translate_off
defparam hex5_obuf_5_.input_async_reset = "none";
defparam hex5_obuf_5_.input_power_up = "low";
defparam hex5_obuf_5_.input_register_mode = "none";
defparam hex5_obuf_5_.input_sync_reset = "none";
defparam hex5_obuf_5_.oe_async_reset = "none";
defparam hex5_obuf_5_.oe_power_up = "low";
defparam hex5_obuf_5_.oe_register_mode = "none";
defparam hex5_obuf_5_.oe_sync_reset = "none";
defparam hex5_obuf_5_.operation_mode = "output";
defparam hex5_obuf_5_.output_async_reset = "none";
defparam hex5_obuf_5_.output_power_up = "low";
defparam hex5_obuf_5_.output_register_mode = "none";
defparam hex5_obuf_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_R3
cycloneii_io hex5_obuf_6_(
	.datain(hex5_dup0_6_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex5[6]));
// synopsys translate_off
defparam hex5_obuf_6_.input_async_reset = "none";
defparam hex5_obuf_6_.input_power_up = "low";
defparam hex5_obuf_6_.input_register_mode = "none";
defparam hex5_obuf_6_.input_sync_reset = "none";
defparam hex5_obuf_6_.oe_async_reset = "none";
defparam hex5_obuf_6_.oe_power_up = "low";
defparam hex5_obuf_6_.oe_register_mode = "none";
defparam hex5_obuf_6_.oe_sync_reset = "none";
defparam hex5_obuf_6_.operation_mode = "output";
defparam hex5_obuf_6_.output_async_reset = "none";
defparam hex5_obuf_6_.output_power_up = "low";
defparam hex5_obuf_6_.output_register_mode = "none";
defparam hex5_obuf_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_R2
cycloneii_io hex6_obuf_0_(
	.datain(hex6_dup0_0_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex6[0]));
// synopsys translate_off
defparam hex6_obuf_0_.input_async_reset = "none";
defparam hex6_obuf_0_.input_power_up = "low";
defparam hex6_obuf_0_.input_register_mode = "none";
defparam hex6_obuf_0_.input_sync_reset = "none";
defparam hex6_obuf_0_.oe_async_reset = "none";
defparam hex6_obuf_0_.oe_power_up = "low";
defparam hex6_obuf_0_.oe_register_mode = "none";
defparam hex6_obuf_0_.oe_sync_reset = "none";
defparam hex6_obuf_0_.operation_mode = "output";
defparam hex6_obuf_0_.output_async_reset = "none";
defparam hex6_obuf_0_.output_power_up = "low";
defparam hex6_obuf_0_.output_register_mode = "none";
defparam hex6_obuf_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P4
cycloneii_io hex6_obuf_1_(
	.datain(hex6_dup0_1_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex6[1]));
// synopsys translate_off
defparam hex6_obuf_1_.input_async_reset = "none";
defparam hex6_obuf_1_.input_power_up = "low";
defparam hex6_obuf_1_.input_register_mode = "none";
defparam hex6_obuf_1_.input_sync_reset = "none";
defparam hex6_obuf_1_.oe_async_reset = "none";
defparam hex6_obuf_1_.oe_power_up = "low";
defparam hex6_obuf_1_.oe_register_mode = "none";
defparam hex6_obuf_1_.oe_sync_reset = "none";
defparam hex6_obuf_1_.operation_mode = "output";
defparam hex6_obuf_1_.output_async_reset = "none";
defparam hex6_obuf_1_.output_power_up = "low";
defparam hex6_obuf_1_.output_register_mode = "none";
defparam hex6_obuf_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P3
cycloneii_io hex6_obuf_2_(
	.datain(hex6_dup0_2_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex6[2]));
// synopsys translate_off
defparam hex6_obuf_2_.input_async_reset = "none";
defparam hex6_obuf_2_.input_power_up = "low";
defparam hex6_obuf_2_.input_register_mode = "none";
defparam hex6_obuf_2_.input_sync_reset = "none";
defparam hex6_obuf_2_.oe_async_reset = "none";
defparam hex6_obuf_2_.oe_power_up = "low";
defparam hex6_obuf_2_.oe_register_mode = "none";
defparam hex6_obuf_2_.oe_sync_reset = "none";
defparam hex6_obuf_2_.operation_mode = "output";
defparam hex6_obuf_2_.output_async_reset = "none";
defparam hex6_obuf_2_.output_power_up = "low";
defparam hex6_obuf_2_.output_register_mode = "none";
defparam hex6_obuf_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_M2
cycloneii_io hex6_obuf_3_(
	.datain(hex6_dup0_3_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex6[3]));
// synopsys translate_off
defparam hex6_obuf_3_.input_async_reset = "none";
defparam hex6_obuf_3_.input_power_up = "low";
defparam hex6_obuf_3_.input_register_mode = "none";
defparam hex6_obuf_3_.input_sync_reset = "none";
defparam hex6_obuf_3_.oe_async_reset = "none";
defparam hex6_obuf_3_.oe_power_up = "low";
defparam hex6_obuf_3_.oe_register_mode = "none";
defparam hex6_obuf_3_.oe_sync_reset = "none";
defparam hex6_obuf_3_.operation_mode = "output";
defparam hex6_obuf_3_.output_async_reset = "none";
defparam hex6_obuf_3_.output_power_up = "low";
defparam hex6_obuf_3_.output_register_mode = "none";
defparam hex6_obuf_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_M3
cycloneii_io hex6_obuf_4_(
	.datain(hex6_dup0_4_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex6[4]));
// synopsys translate_off
defparam hex6_obuf_4_.input_async_reset = "none";
defparam hex6_obuf_4_.input_power_up = "low";
defparam hex6_obuf_4_.input_register_mode = "none";
defparam hex6_obuf_4_.input_sync_reset = "none";
defparam hex6_obuf_4_.oe_async_reset = "none";
defparam hex6_obuf_4_.oe_power_up = "low";
defparam hex6_obuf_4_.oe_register_mode = "none";
defparam hex6_obuf_4_.oe_sync_reset = "none";
defparam hex6_obuf_4_.operation_mode = "output";
defparam hex6_obuf_4_.output_async_reset = "none";
defparam hex6_obuf_4_.output_power_up = "low";
defparam hex6_obuf_4_.output_register_mode = "none";
defparam hex6_obuf_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_M5
cycloneii_io hex6_obuf_5_(
	.datain(hex6_dup0_5_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex6[5]));
// synopsys translate_off
defparam hex6_obuf_5_.input_async_reset = "none";
defparam hex6_obuf_5_.input_power_up = "low";
defparam hex6_obuf_5_.input_register_mode = "none";
defparam hex6_obuf_5_.input_sync_reset = "none";
defparam hex6_obuf_5_.oe_async_reset = "none";
defparam hex6_obuf_5_.oe_power_up = "low";
defparam hex6_obuf_5_.oe_register_mode = "none";
defparam hex6_obuf_5_.oe_sync_reset = "none";
defparam hex6_obuf_5_.operation_mode = "output";
defparam hex6_obuf_5_.output_async_reset = "none";
defparam hex6_obuf_5_.output_power_up = "low";
defparam hex6_obuf_5_.output_register_mode = "none";
defparam hex6_obuf_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_M4
cycloneii_io hex6_obuf_6_(
	.datain(hex6_dup0_6_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex6[6]));
// synopsys translate_off
defparam hex6_obuf_6_.input_async_reset = "none";
defparam hex6_obuf_6_.input_power_up = "low";
defparam hex6_obuf_6_.input_register_mode = "none";
defparam hex6_obuf_6_.input_sync_reset = "none";
defparam hex6_obuf_6_.oe_async_reset = "none";
defparam hex6_obuf_6_.oe_power_up = "low";
defparam hex6_obuf_6_.oe_register_mode = "none";
defparam hex6_obuf_6_.oe_sync_reset = "none";
defparam hex6_obuf_6_.operation_mode = "output";
defparam hex6_obuf_6_.output_async_reset = "none";
defparam hex6_obuf_6_.output_power_up = "low";
defparam hex6_obuf_6_.output_register_mode = "none";
defparam hex6_obuf_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_L3
cycloneii_io hex7_obuf_0_(
	.datain(hex7_dup0_0_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex7[0]));
// synopsys translate_off
defparam hex7_obuf_0_.input_async_reset = "none";
defparam hex7_obuf_0_.input_power_up = "low";
defparam hex7_obuf_0_.input_register_mode = "none";
defparam hex7_obuf_0_.input_sync_reset = "none";
defparam hex7_obuf_0_.oe_async_reset = "none";
defparam hex7_obuf_0_.oe_power_up = "low";
defparam hex7_obuf_0_.oe_register_mode = "none";
defparam hex7_obuf_0_.oe_sync_reset = "none";
defparam hex7_obuf_0_.operation_mode = "output";
defparam hex7_obuf_0_.output_async_reset = "none";
defparam hex7_obuf_0_.output_power_up = "low";
defparam hex7_obuf_0_.output_register_mode = "none";
defparam hex7_obuf_0_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_L2
cycloneii_io hex7_obuf_1_(
	.datain(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex7[1]));
// synopsys translate_off
defparam hex7_obuf_1_.input_async_reset = "none";
defparam hex7_obuf_1_.input_power_up = "low";
defparam hex7_obuf_1_.input_register_mode = "none";
defparam hex7_obuf_1_.input_sync_reset = "none";
defparam hex7_obuf_1_.oe_async_reset = "none";
defparam hex7_obuf_1_.oe_power_up = "low";
defparam hex7_obuf_1_.oe_register_mode = "none";
defparam hex7_obuf_1_.oe_sync_reset = "none";
defparam hex7_obuf_1_.operation_mode = "output";
defparam hex7_obuf_1_.output_async_reset = "none";
defparam hex7_obuf_1_.output_power_up = "low";
defparam hex7_obuf_1_.output_register_mode = "none";
defparam hex7_obuf_1_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_L9
cycloneii_io hex7_obuf_2_(
	.datain(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex7[2]));
// synopsys translate_off
defparam hex7_obuf_2_.input_async_reset = "none";
defparam hex7_obuf_2_.input_power_up = "low";
defparam hex7_obuf_2_.input_register_mode = "none";
defparam hex7_obuf_2_.input_sync_reset = "none";
defparam hex7_obuf_2_.oe_async_reset = "none";
defparam hex7_obuf_2_.oe_power_up = "low";
defparam hex7_obuf_2_.oe_register_mode = "none";
defparam hex7_obuf_2_.oe_sync_reset = "none";
defparam hex7_obuf_2_.operation_mode = "output";
defparam hex7_obuf_2_.output_async_reset = "none";
defparam hex7_obuf_2_.output_power_up = "low";
defparam hex7_obuf_2_.output_register_mode = "none";
defparam hex7_obuf_2_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_L6
cycloneii_io hex7_obuf_3_(
	.datain(hex7_dup0_0_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex7[3]));
// synopsys translate_off
defparam hex7_obuf_3_.input_async_reset = "none";
defparam hex7_obuf_3_.input_power_up = "low";
defparam hex7_obuf_3_.input_register_mode = "none";
defparam hex7_obuf_3_.input_sync_reset = "none";
defparam hex7_obuf_3_.oe_async_reset = "none";
defparam hex7_obuf_3_.oe_power_up = "low";
defparam hex7_obuf_3_.oe_register_mode = "none";
defparam hex7_obuf_3_.oe_sync_reset = "none";
defparam hex7_obuf_3_.operation_mode = "output";
defparam hex7_obuf_3_.output_async_reset = "none";
defparam hex7_obuf_3_.output_power_up = "low";
defparam hex7_obuf_3_.output_register_mode = "none";
defparam hex7_obuf_3_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_L7
cycloneii_io hex7_obuf_4_(
	.datain(hex7_dup0_0_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex7[4]));
// synopsys translate_off
defparam hex7_obuf_4_.input_async_reset = "none";
defparam hex7_obuf_4_.input_power_up = "low";
defparam hex7_obuf_4_.input_register_mode = "none";
defparam hex7_obuf_4_.input_sync_reset = "none";
defparam hex7_obuf_4_.oe_async_reset = "none";
defparam hex7_obuf_4_.oe_power_up = "low";
defparam hex7_obuf_4_.oe_register_mode = "none";
defparam hex7_obuf_4_.oe_sync_reset = "none";
defparam hex7_obuf_4_.operation_mode = "output";
defparam hex7_obuf_4_.output_async_reset = "none";
defparam hex7_obuf_4_.output_power_up = "low";
defparam hex7_obuf_4_.output_register_mode = "none";
defparam hex7_obuf_4_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P9
cycloneii_io hex7_obuf_5_(
	.datain(hex7_dup0_0_),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex7[5]));
// synopsys translate_off
defparam hex7_obuf_5_.input_async_reset = "none";
defparam hex7_obuf_5_.input_power_up = "low";
defparam hex7_obuf_5_.input_register_mode = "none";
defparam hex7_obuf_5_.input_sync_reset = "none";
defparam hex7_obuf_5_.oe_async_reset = "none";
defparam hex7_obuf_5_.oe_power_up = "low";
defparam hex7_obuf_5_.oe_register_mode = "none";
defparam hex7_obuf_5_.oe_sync_reset = "none";
defparam hex7_obuf_5_.operation_mode = "output";
defparam hex7_obuf_5_.output_async_reset = "none";
defparam hex7_obuf_5_.output_power_up = "low";
defparam hex7_obuf_5_.output_register_mode = "none";
defparam hex7_obuf_5_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_N9
cycloneii_io hex7_obuf_6_(
	.datain(vcc),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(hex7[6]));
// synopsys translate_off
defparam hex7_obuf_6_.input_async_reset = "none";
defparam hex7_obuf_6_.input_power_up = "low";
defparam hex7_obuf_6_.input_register_mode = "none";
defparam hex7_obuf_6_.input_sync_reset = "none";
defparam hex7_obuf_6_.oe_async_reset = "none";
defparam hex7_obuf_6_.oe_power_up = "low";
defparam hex7_obuf_6_.oe_register_mode = "none";
defparam hex7_obuf_6_.oe_sync_reset = "none";
defparam hex7_obuf_6_.operation_mode = "output";
defparam hex7_obuf_6_.output_async_reset = "none";
defparam hex7_obuf_6_.output_power_up = "low";
defparam hex7_obuf_6_.output_register_mode = "none";
defparam hex7_obuf_6_.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_A5
cycloneii_io aud_xck_obuf(
	.datain(\u_audio_dac_p1_altpll|_clk1~clkctrl_outclk ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(aud_xck));
// synopsys translate_off
defparam aud_xck_obuf.input_async_reset = "none";
defparam aud_xck_obuf.input_power_up = "low";
defparam aud_xck_obuf.input_register_mode = "none";
defparam aud_xck_obuf.input_sync_reset = "none";
defparam aud_xck_obuf.oe_async_reset = "none";
defparam aud_xck_obuf.oe_power_up = "low";
defparam aud_xck_obuf.oe_register_mode = "none";
defparam aud_xck_obuf.oe_sync_reset = "none";
defparam aud_xck_obuf.operation_mode = "output";
defparam aud_xck_obuf.output_async_reset = "none";
defparam aud_xck_obuf.output_power_up = "low";
defparam aud_xck_obuf.output_register_mode = "none";
defparam aud_xck_obuf.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_A4
cycloneii_io aud_dacdat_obuf(
	.datain(aud_dacdat_dup0),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(aud_dacdat));
// synopsys translate_off
defparam aud_dacdat_obuf.input_async_reset = "none";
defparam aud_dacdat_obuf.input_power_up = "low";
defparam aud_dacdat_obuf.input_register_mode = "none";
defparam aud_dacdat_obuf.input_sync_reset = "none";
defparam aud_dacdat_obuf.oe_async_reset = "none";
defparam aud_dacdat_obuf.oe_power_up = "low";
defparam aud_dacdat_obuf.oe_register_mode = "none";
defparam aud_dacdat_obuf.oe_sync_reset = "none";
defparam aud_dacdat_obuf.operation_mode = "output";
defparam aud_dacdat_obuf.output_async_reset = "none";
defparam aud_dacdat_obuf.output_power_up = "low";
defparam aud_dacdat_obuf.output_register_mode = "none";
defparam aud_dacdat_obuf.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_C6
cycloneii_io aud_daclrck_obuf(
	.datain(aud_adclrck_dup0),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(aud_daclrck));
// synopsys translate_off
defparam aud_daclrck_obuf.input_async_reset = "none";
defparam aud_daclrck_obuf.input_power_up = "low";
defparam aud_daclrck_obuf.input_register_mode = "none";
defparam aud_daclrck_obuf.input_sync_reset = "none";
defparam aud_daclrck_obuf.oe_async_reset = "none";
defparam aud_daclrck_obuf.oe_power_up = "low";
defparam aud_daclrck_obuf.oe_register_mode = "none";
defparam aud_daclrck_obuf.oe_sync_reset = "none";
defparam aud_daclrck_obuf.operation_mode = "output";
defparam aud_daclrck_obuf.output_async_reset = "none";
defparam aud_daclrck_obuf.output_power_up = "low";
defparam aud_daclrck_obuf.output_register_mode = "none";
defparam aud_daclrck_obuf.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_C5
cycloneii_io aud_adclrck_obuf(
	.datain(aud_adclrck_dup0),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(aud_adclrck));
// synopsys translate_off
defparam aud_adclrck_obuf.input_async_reset = "none";
defparam aud_adclrck_obuf.input_power_up = "low";
defparam aud_adclrck_obuf.input_register_mode = "none";
defparam aud_adclrck_obuf.input_sync_reset = "none";
defparam aud_adclrck_obuf.oe_async_reset = "none";
defparam aud_adclrck_obuf.oe_power_up = "low";
defparam aud_adclrck_obuf.oe_register_mode = "none";
defparam aud_adclrck_obuf.oe_sync_reset = "none";
defparam aud_adclrck_obuf.operation_mode = "output";
defparam aud_adclrck_obuf.output_async_reset = "none";
defparam aud_adclrck_obuf.output_power_up = "low";
defparam aud_adclrck_obuf.output_register_mode = "none";
defparam aud_adclrck_obuf.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_A6
cycloneii_io i2c_sclk_obuf(
	.datain(\u_i2c_av_config|u0|p_i2c_sclk ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(i2c_sclk));
// synopsys translate_off
defparam i2c_sclk_obuf.input_async_reset = "none";
defparam i2c_sclk_obuf.input_power_up = "low";
defparam i2c_sclk_obuf.input_register_mode = "none";
defparam i2c_sclk_obuf.input_sync_reset = "none";
defparam i2c_sclk_obuf.oe_async_reset = "none";
defparam i2c_sclk_obuf.oe_power_up = "low";
defparam i2c_sclk_obuf.oe_register_mode = "none";
defparam i2c_sclk_obuf.oe_sync_reset = "none";
defparam i2c_sclk_obuf.operation_mode = "output";
defparam i2c_sclk_obuf.output_async_reset = "none";
defparam i2c_sclk_obuf.output_power_up = "low";
defparam i2c_sclk_obuf.output_register_mode = "none";
defparam i2c_sclk_obuf.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_B6
cycloneii_io u_i2c_av_config_u0_ix31977z43919(
	.datain(!\u_i2c_av_config|u0|nx51857z1 ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(i2c_sdat));
// synopsys translate_off
defparam u_i2c_av_config_u0_ix31977z43919.input_async_reset = "none";
defparam u_i2c_av_config_u0_ix31977z43919.input_power_up = "low";
defparam u_i2c_av_config_u0_ix31977z43919.input_register_mode = "none";
defparam u_i2c_av_config_u0_ix31977z43919.input_sync_reset = "none";
defparam u_i2c_av_config_u0_ix31977z43919.oe_async_reset = "none";
defparam u_i2c_av_config_u0_ix31977z43919.oe_power_up = "low";
defparam u_i2c_av_config_u0_ix31977z43919.oe_register_mode = "none";
defparam u_i2c_av_config_u0_ix31977z43919.oe_sync_reset = "none";
defparam u_i2c_av_config_u0_ix31977z43919.open_drain_output = "true";
defparam u_i2c_av_config_u0_ix31977z43919.operation_mode = "bidir";
defparam u_i2c_av_config_u0_ix31977z43919.output_async_reset = "none";
defparam u_i2c_av_config_u0_ix31977z43919.output_power_up = "low";
defparam u_i2c_av_config_u0_ix31977z43919.output_register_mode = "none";
defparam u_i2c_av_config_u0_ix31977z43919.output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_B4
cycloneii_io \aud_bclk~I (
	.datain(aud_bclk_dup0),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(aud_bclk));
// synopsys translate_off
defparam \aud_bclk~I .input_async_reset = "none";
defparam \aud_bclk~I .input_power_up = "low";
defparam \aud_bclk~I .input_register_mode = "none";
defparam \aud_bclk~I .input_sync_reset = "none";
defparam \aud_bclk~I .oe_async_reset = "none";
defparam \aud_bclk~I .oe_power_up = "low";
defparam \aud_bclk~I .oe_register_mode = "none";
defparam \aud_bclk~I .oe_sync_reset = "none";
defparam \aud_bclk~I .operation_mode = "bidir";
defparam \aud_bclk~I .output_async_reset = "none";
defparam \aud_bclk~I .output_power_up = "low";
defparam \aud_bclk~I .output_register_mode = "none";
defparam \aud_bclk~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_N2
cycloneii_io \clock_50~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(clock_50));
// synopsys translate_off
defparam \clock_50~I .input_async_reset = "none";
defparam \clock_50~I .input_power_up = "low";
defparam \clock_50~I .input_register_mode = "none";
defparam \clock_50~I .input_sync_reset = "none";
defparam \clock_50~I .oe_async_reset = "none";
defparam \clock_50~I .oe_power_up = "low";
defparam \clock_50~I .oe_register_mode = "none";
defparam \clock_50~I .oe_sync_reset = "none";
defparam \clock_50~I .operation_mode = "input";
defparam \clock_50~I .output_async_reset = "none";
defparam \clock_50~I .output_power_up = "low";
defparam \clock_50~I .output_register_mode = "none";
defparam \clock_50~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_N23
cycloneii_io \key[1]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(key[1]));
// synopsys translate_off
defparam \key[1]~I .input_async_reset = "none";
defparam \key[1]~I .input_power_up = "low";
defparam \key[1]~I .input_register_mode = "none";
defparam \key[1]~I .input_sync_reset = "none";
defparam \key[1]~I .oe_async_reset = "none";
defparam \key[1]~I .oe_power_up = "low";
defparam \key[1]~I .oe_register_mode = "none";
defparam \key[1]~I .oe_sync_reset = "none";
defparam \key[1]~I .operation_mode = "input";
defparam \key[1]~I .output_async_reset = "none";
defparam \key[1]~I .output_power_up = "low";
defparam \key[1]~I .output_register_mode = "none";
defparam \key[1]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P23
cycloneii_io \key[2]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(key[2]));
// synopsys translate_off
defparam \key[2]~I .input_async_reset = "none";
defparam \key[2]~I .input_power_up = "low";
defparam \key[2]~I .input_register_mode = "none";
defparam \key[2]~I .input_sync_reset = "none";
defparam \key[2]~I .oe_async_reset = "none";
defparam \key[2]~I .oe_power_up = "low";
defparam \key[2]~I .oe_register_mode = "none";
defparam \key[2]~I .oe_sync_reset = "none";
defparam \key[2]~I .operation_mode = "input";
defparam \key[2]~I .output_async_reset = "none";
defparam \key[2]~I .output_power_up = "low";
defparam \key[2]~I .output_register_mode = "none";
defparam \key[2]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_W26
cycloneii_io \key[3]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(key[3]));
// synopsys translate_off
defparam \key[3]~I .input_async_reset = "none";
defparam \key[3]~I .input_power_up = "low";
defparam \key[3]~I .input_register_mode = "none";
defparam \key[3]~I .input_sync_reset = "none";
defparam \key[3]~I .oe_async_reset = "none";
defparam \key[3]~I .oe_power_up = "low";
defparam \key[3]~I .oe_register_mode = "none";
defparam \key[3]~I .oe_sync_reset = "none";
defparam \key[3]~I .operation_mode = "input";
defparam \key[3]~I .output_async_reset = "none";
defparam \key[3]~I .output_power_up = "low";
defparam \key[3]~I .output_register_mode = "none";
defparam \key[3]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_C13
cycloneii_io \sw[7]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[7]));
// synopsys translate_off
defparam \sw[7]~I .input_async_reset = "none";
defparam \sw[7]~I .input_power_up = "low";
defparam \sw[7]~I .input_register_mode = "none";
defparam \sw[7]~I .input_sync_reset = "none";
defparam \sw[7]~I .oe_async_reset = "none";
defparam \sw[7]~I .oe_power_up = "low";
defparam \sw[7]~I .oe_register_mode = "none";
defparam \sw[7]~I .oe_sync_reset = "none";
defparam \sw[7]~I .operation_mode = "input";
defparam \sw[7]~I .output_async_reset = "none";
defparam \sw[7]~I .output_power_up = "low";
defparam \sw[7]~I .output_register_mode = "none";
defparam \sw[7]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_B13
cycloneii_io \sw[8]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[8]));
// synopsys translate_off
defparam \sw[8]~I .input_async_reset = "none";
defparam \sw[8]~I .input_power_up = "low";
defparam \sw[8]~I .input_register_mode = "none";
defparam \sw[8]~I .input_sync_reset = "none";
defparam \sw[8]~I .oe_async_reset = "none";
defparam \sw[8]~I .oe_power_up = "low";
defparam \sw[8]~I .oe_register_mode = "none";
defparam \sw[8]~I .oe_sync_reset = "none";
defparam \sw[8]~I .operation_mode = "input";
defparam \sw[8]~I .output_async_reset = "none";
defparam \sw[8]~I .output_power_up = "low";
defparam \sw[8]~I .output_register_mode = "none";
defparam \sw[8]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_A13
cycloneii_io \sw[9]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[9]));
// synopsys translate_off
defparam \sw[9]~I .input_async_reset = "none";
defparam \sw[9]~I .input_power_up = "low";
defparam \sw[9]~I .input_register_mode = "none";
defparam \sw[9]~I .input_sync_reset = "none";
defparam \sw[9]~I .oe_async_reset = "none";
defparam \sw[9]~I .oe_power_up = "low";
defparam \sw[9]~I .oe_register_mode = "none";
defparam \sw[9]~I .oe_sync_reset = "none";
defparam \sw[9]~I .operation_mode = "input";
defparam \sw[9]~I .output_async_reset = "none";
defparam \sw[9]~I .output_power_up = "low";
defparam \sw[9]~I .output_register_mode = "none";
defparam \sw[9]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_N1
cycloneii_io \sw[10]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[10]));
// synopsys translate_off
defparam \sw[10]~I .input_async_reset = "none";
defparam \sw[10]~I .input_power_up = "low";
defparam \sw[10]~I .input_register_mode = "none";
defparam \sw[10]~I .input_sync_reset = "none";
defparam \sw[10]~I .oe_async_reset = "none";
defparam \sw[10]~I .oe_power_up = "low";
defparam \sw[10]~I .oe_register_mode = "none";
defparam \sw[10]~I .oe_sync_reset = "none";
defparam \sw[10]~I .operation_mode = "input";
defparam \sw[10]~I .output_async_reset = "none";
defparam \sw[10]~I .output_power_up = "low";
defparam \sw[10]~I .output_register_mode = "none";
defparam \sw[10]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P1
cycloneii_io \sw[11]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[11]));
// synopsys translate_off
defparam \sw[11]~I .input_async_reset = "none";
defparam \sw[11]~I .input_power_up = "low";
defparam \sw[11]~I .input_register_mode = "none";
defparam \sw[11]~I .input_sync_reset = "none";
defparam \sw[11]~I .oe_async_reset = "none";
defparam \sw[11]~I .oe_power_up = "low";
defparam \sw[11]~I .oe_register_mode = "none";
defparam \sw[11]~I .oe_sync_reset = "none";
defparam \sw[11]~I .operation_mode = "input";
defparam \sw[11]~I .output_async_reset = "none";
defparam \sw[11]~I .output_power_up = "low";
defparam \sw[11]~I .output_register_mode = "none";
defparam \sw[11]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_P2
cycloneii_io \sw[12]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[12]));
// synopsys translate_off
defparam \sw[12]~I .input_async_reset = "none";
defparam \sw[12]~I .input_power_up = "low";
defparam \sw[12]~I .input_register_mode = "none";
defparam \sw[12]~I .input_sync_reset = "none";
defparam \sw[12]~I .oe_async_reset = "none";
defparam \sw[12]~I .oe_power_up = "low";
defparam \sw[12]~I .oe_register_mode = "none";
defparam \sw[12]~I .oe_sync_reset = "none";
defparam \sw[12]~I .operation_mode = "input";
defparam \sw[12]~I .output_async_reset = "none";
defparam \sw[12]~I .output_power_up = "low";
defparam \sw[12]~I .output_register_mode = "none";
defparam \sw[12]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_T7
cycloneii_io \sw[13]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[13]));
// synopsys translate_off
defparam \sw[13]~I .input_async_reset = "none";
defparam \sw[13]~I .input_power_up = "low";
defparam \sw[13]~I .input_register_mode = "none";
defparam \sw[13]~I .input_sync_reset = "none";
defparam \sw[13]~I .oe_async_reset = "none";
defparam \sw[13]~I .oe_power_up = "low";
defparam \sw[13]~I .oe_register_mode = "none";
defparam \sw[13]~I .oe_sync_reset = "none";
defparam \sw[13]~I .operation_mode = "input";
defparam \sw[13]~I .output_async_reset = "none";
defparam \sw[13]~I .output_power_up = "low";
defparam \sw[13]~I .output_register_mode = "none";
defparam \sw[13]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_U3
cycloneii_io \sw[14]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[14]));
// synopsys translate_off
defparam \sw[14]~I .input_async_reset = "none";
defparam \sw[14]~I .input_power_up = "low";
defparam \sw[14]~I .input_register_mode = "none";
defparam \sw[14]~I .input_sync_reset = "none";
defparam \sw[14]~I .oe_async_reset = "none";
defparam \sw[14]~I .oe_power_up = "low";
defparam \sw[14]~I .oe_register_mode = "none";
defparam \sw[14]~I .oe_sync_reset = "none";
defparam \sw[14]~I .operation_mode = "input";
defparam \sw[14]~I .output_async_reset = "none";
defparam \sw[14]~I .output_power_up = "low";
defparam \sw[14]~I .output_register_mode = "none";
defparam \sw[14]~I .output_sync_reset = "none";
// synopsys translate_on

// atom is at PIN_U4
cycloneii_io \sw[15]~I (
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.differentialin(gnd),
	.linkin(gnd),
	.devclrn(devclrn),
	.devpor(devpor),
	.devoe(devoe),
	.combout(),
	.regout(),
	.differentialout(),
	.linkout(),
	.padio(sw[15]));
// synopsys translate_off
defparam \sw[15]~I .input_async_reset = "none";
defparam \sw[15]~I .input_power_up = "low";
defparam \sw[15]~I .input_register_mode = "none";
defparam \sw[15]~I .input_sync_reset = "none";
defparam \sw[15]~I .oe_async_reset = "none";
defparam \sw[15]~I .oe_power_up = "low";
defparam \sw[15]~I .oe_register_mode = "none";
defparam \sw[15]~I .oe_sync_reset = "none";
defparam \sw[15]~I .operation_mode = "input";
defparam \sw[15]~I .output_async_reset = "none";
defparam \sw[15]~I .output_power_up = "low";
defparam \sw[15]~I .output_register_mode = "none";
defparam \sw[15]~I .output_sync_reset = "none";
// synopsys translate_on

endmodule
